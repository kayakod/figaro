magic
tech sky130A
magscale 1 2
timestamp 1654677594
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 309134 700884 309140 700936
rect 309192 700924 309198 700936
rect 364978 700924 364984 700936
rect 309192 700896 364984 700924
rect 309192 700884 309198 700896
rect 364978 700884 364984 700896
rect 365036 700884 365042 700936
rect 313274 700816 313280 700868
rect 313332 700856 313338 700868
rect 397454 700856 397460 700868
rect 313332 700828 397460 700856
rect 313332 700816 313338 700828
rect 397454 700816 397460 700828
rect 397512 700816 397518 700868
rect 317414 700748 317420 700800
rect 317472 700788 317478 700800
rect 413646 700788 413652 700800
rect 317472 700760 413652 700788
rect 317472 700748 317478 700760
rect 413646 700748 413652 700760
rect 413704 700748 413710 700800
rect 322934 700680 322940 700732
rect 322992 700720 322998 700732
rect 429838 700720 429844 700732
rect 322992 700692 429844 700720
rect 322992 700680 322998 700692
rect 429838 700680 429844 700692
rect 429896 700680 429902 700732
rect 327074 700612 327080 700664
rect 327132 700652 327138 700664
rect 462314 700652 462320 700664
rect 327132 700624 462320 700652
rect 327132 700612 327138 700624
rect 462314 700612 462320 700624
rect 462372 700612 462378 700664
rect 331306 700544 331312 700596
rect 331364 700584 331370 700596
rect 478506 700584 478512 700596
rect 331364 700556 478512 700584
rect 331364 700544 331370 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 335354 700476 335360 700528
rect 335412 700516 335418 700528
rect 494790 700516 494796 700528
rect 335412 700488 494796 700516
rect 335412 700476 335418 700488
rect 494790 700476 494796 700488
rect 494848 700476 494854 700528
rect 340874 700408 340880 700460
rect 340932 700448 340938 700460
rect 527174 700448 527180 700460
rect 340932 700420 527180 700448
rect 340932 700408 340938 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 300854 700340 300860 700392
rect 300912 700380 300918 700392
rect 332502 700380 332508 700392
rect 300912 700352 332508 700380
rect 300912 700340 300918 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 345014 700340 345020 700392
rect 345072 700380 345078 700392
rect 543458 700380 543464 700392
rect 345072 700352 543464 700380
rect 345072 700340 345078 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 279418 700312 279424 700324
rect 267700 700284 279424 700312
rect 267700 700272 267706 700284
rect 279418 700272 279424 700284
rect 279476 700272 279482 700324
rect 295334 700272 295340 700324
rect 295392 700312 295398 700324
rect 300118 700312 300124 700324
rect 295392 700284 300124 700312
rect 295392 700272 295398 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 304994 700272 305000 700324
rect 305052 700312 305058 700324
rect 348786 700312 348792 700324
rect 305052 700284 348792 700312
rect 305052 700272 305058 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 349154 700272 349160 700324
rect 349212 700312 349218 700324
rect 559650 700312 559656 700324
rect 349212 700284 559656 700312
rect 349212 700272 349218 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 353938 683136 353944 683188
rect 353996 683176 354002 683188
rect 579614 683176 579620 683188
rect 353996 683148 579620 683176
rect 353996 683136 354002 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 360838 670692 360844 670744
rect 360896 670732 360902 670744
rect 580166 670732 580172 670744
rect 360896 670704 580172 670732
rect 360896 670692 360902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 367738 643084 367744 643136
rect 367796 643124 367802 643136
rect 580166 643124 580172 643136
rect 367796 643096 580172 643124
rect 367796 643084 367802 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3326 632068 3332 632120
rect 3384 632108 3390 632120
rect 32398 632108 32404 632120
rect 3384 632080 32404 632108
rect 3384 632068 3390 632080
rect 32398 632068 32404 632080
rect 32456 632068 32462 632120
rect 374638 630640 374644 630692
rect 374696 630680 374702 630692
rect 579982 630680 579988 630692
rect 374696 630652 579988 630680
rect 374696 630640 374702 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3326 618264 3332 618316
rect 3384 618304 3390 618316
rect 22738 618304 22744 618316
rect 3384 618276 22744 618304
rect 3384 618264 3390 618276
rect 22738 618264 22744 618276
rect 22796 618264 22802 618316
rect 381538 616836 381544 616888
rect 381596 616876 381602 616888
rect 580166 616876 580172 616888
rect 381596 616848 580172 616876
rect 381596 616836 381602 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 14458 605860 14464 605872
rect 3384 605832 14464 605860
rect 3384 605820 3390 605832
rect 14458 605820 14464 605832
rect 14516 605820 14522 605872
rect 3142 579776 3148 579828
rect 3200 579816 3206 579828
rect 7558 579816 7564 579828
rect 3200 579788 7564 579816
rect 3200 579776 3206 579788
rect 7558 579776 7564 579788
rect 7616 579776 7622 579828
rect 359458 563048 359464 563100
rect 359516 563088 359522 563100
rect 580166 563088 580172 563100
rect 359516 563060 580172 563088
rect 359516 563048 359522 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 364978 536800 364984 536852
rect 365036 536840 365042 536852
rect 580166 536840 580172 536852
rect 365036 536812 580172 536840
rect 365036 536800 365042 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 43438 527184 43444 527196
rect 3016 527156 43444 527184
rect 3016 527144 3022 527156
rect 43438 527144 43444 527156
rect 43496 527144 43502 527196
rect 373258 524424 373264 524476
rect 373316 524464 373322 524476
rect 580166 524464 580172 524476
rect 373316 524436 580172 524464
rect 373316 524424 373322 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 25498 514808 25504 514820
rect 3384 514780 25504 514808
rect 3384 514768 3390 514780
rect 25498 514768 25504 514780
rect 25556 514768 25562 514820
rect 356698 510620 356704 510672
rect 356756 510660 356762 510672
rect 580166 510660 580172 510672
rect 356756 510632 580172 510660
rect 356756 510620 356762 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 17218 501004 17224 501016
rect 3292 500976 17224 501004
rect 3292 500964 3298 500976
rect 17218 500964 17224 500976
rect 17276 500964 17282 501016
rect 3326 475192 3332 475244
rect 3384 475232 3390 475244
rect 8938 475232 8944 475244
rect 3384 475204 8944 475232
rect 3384 475192 3390 475204
rect 8938 475192 8944 475204
rect 8996 475192 9002 475244
rect 355318 456764 355324 456816
rect 355376 456804 355382 456816
rect 580166 456804 580172 456816
rect 355376 456776 580172 456804
rect 355376 456764 355382 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 371878 430584 371884 430636
rect 371936 430624 371942 430636
rect 580166 430624 580172 430636
rect 371936 430596 580172 430624
rect 371936 430584 371942 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 31018 422328 31024 422340
rect 3016 422300 31024 422328
rect 3016 422288 3022 422300
rect 31018 422288 31024 422300
rect 31076 422288 31082 422340
rect 378778 418140 378784 418192
rect 378836 418180 378842 418192
rect 580166 418180 580172 418192
rect 378836 418152 580172 418180
rect 378836 418140 378842 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 26878 409884 26884 409896
rect 3384 409856 26884 409884
rect 3384 409844 3390 409856
rect 26878 409844 26884 409856
rect 26936 409844 26942 409896
rect 363598 404336 363604 404388
rect 363656 404376 363662 404388
rect 580166 404376 580172 404388
rect 363656 404348 580172 404376
rect 363656 404336 363662 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 18598 397508 18604 397520
rect 3384 397480 18604 397508
rect 3384 397468 3390 397480
rect 18598 397468 18604 397480
rect 18656 397468 18662 397520
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 10318 371260 10324 371272
rect 3384 371232 10324 371260
rect 3384 371220 3390 371232
rect 10318 371220 10324 371232
rect 10376 371220 10382 371272
rect 354030 364352 354036 364404
rect 354088 364392 354094 364404
rect 580166 364392 580172 364404
rect 354088 364364 580172 364392
rect 354088 364352 354094 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 369118 324300 369124 324352
rect 369176 324340 369182 324352
rect 579982 324340 579988 324352
rect 369176 324312 579988 324340
rect 369176 324300 369182 324312
rect 579982 324300 579988 324312
rect 580040 324300 580046 324352
rect 3142 318792 3148 318844
rect 3200 318832 3206 318844
rect 221458 318832 221464 318844
rect 3200 318804 221464 318832
rect 3200 318792 3206 318804
rect 221458 318792 221464 318804
rect 221516 318792 221522 318844
rect 377398 311856 377404 311908
rect 377456 311896 377462 311908
rect 579798 311896 579804 311908
rect 377456 311868 579804 311896
rect 377456 311856 377462 311868
rect 579798 311856 579804 311868
rect 579856 311856 579862 311908
rect 3326 304988 3332 305040
rect 3384 305028 3390 305040
rect 28258 305028 28264 305040
rect 3384 305000 28264 305028
rect 3384 304988 3390 305000
rect 28258 304988 28264 305000
rect 28316 304988 28322 305040
rect 442258 298120 442264 298172
rect 442316 298160 442322 298172
rect 580166 298160 580172 298172
rect 442316 298132 580172 298160
rect 442316 298120 442322 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 21358 292584 21364 292596
rect 3384 292556 21364 292584
rect 3384 292544 3390 292556
rect 21358 292544 21364 292556
rect 21416 292544 21422 292596
rect 3234 266364 3240 266416
rect 3292 266404 3298 266416
rect 13078 266404 13084 266416
rect 3292 266376 13084 266404
rect 3292 266364 3298 266376
rect 13078 266364 13084 266376
rect 13136 266364 13142 266416
rect 218054 263508 218060 263560
rect 218112 263548 218118 263560
rect 278590 263548 278596 263560
rect 218112 263520 278596 263548
rect 218112 263508 218118 263520
rect 278590 263508 278596 263520
rect 278648 263508 278654 263560
rect 201494 263440 201500 263492
rect 201552 263480 201558 263492
rect 274174 263480 274180 263492
rect 201552 263452 274180 263480
rect 201552 263440 201558 263452
rect 274174 263440 274180 263452
rect 274232 263440 274238 263492
rect 169754 263372 169760 263424
rect 169812 263412 169818 263424
rect 269758 263412 269764 263424
rect 169812 263384 269764 263412
rect 169812 263372 169818 263384
rect 269758 263372 269764 263384
rect 269816 263372 269822 263424
rect 153194 263304 153200 263356
rect 153252 263344 153258 263356
rect 265342 263344 265348 263356
rect 153252 263316 265348 263344
rect 153252 263304 153258 263316
rect 265342 263304 265348 263316
rect 265400 263304 265406 263356
rect 136634 263236 136640 263288
rect 136692 263276 136698 263288
rect 260834 263276 260840 263288
rect 136692 263248 260840 263276
rect 136692 263236 136698 263248
rect 260834 263236 260840 263248
rect 260892 263236 260898 263288
rect 104894 263168 104900 263220
rect 104952 263208 104958 263220
rect 256418 263208 256424 263220
rect 104952 263180 256424 263208
rect 104952 263168 104958 263180
rect 256418 263168 256424 263180
rect 256476 263168 256482 263220
rect 88334 263100 88340 263152
rect 88392 263140 88398 263152
rect 252002 263140 252008 263152
rect 88392 263112 252008 263140
rect 88392 263100 88398 263112
rect 252002 263100 252008 263112
rect 252060 263100 252066 263152
rect 71774 263032 71780 263084
rect 71832 263072 71838 263084
rect 247494 263072 247500 263084
rect 71832 263044 247500 263072
rect 71832 263032 71838 263044
rect 247494 263032 247500 263044
rect 247552 263032 247558 263084
rect 40034 262964 40040 263016
rect 40092 263004 40098 263016
rect 243078 263004 243084 263016
rect 40092 262976 243084 263004
rect 40092 262964 40098 262976
rect 243078 262964 243084 262976
rect 243136 262964 243142 263016
rect 282914 262964 282920 263016
rect 282972 263004 282978 263016
rect 291930 263004 291936 263016
rect 282972 262976 291936 263004
rect 282972 262964 282978 262976
rect 291930 262964 291936 262976
rect 291988 262964 291994 263016
rect 23474 262896 23480 262948
rect 23532 262936 23538 262948
rect 238662 262936 238668 262948
rect 23532 262908 238668 262936
rect 23532 262896 23538 262908
rect 238662 262896 238668 262908
rect 238720 262896 238726 262948
rect 279418 262896 279424 262948
rect 279476 262936 279482 262948
rect 287514 262936 287520 262948
rect 279476 262908 287520 262936
rect 279476 262896 279482 262908
rect 287514 262896 287520 262908
rect 287572 262896 287578 262948
rect 6914 262828 6920 262880
rect 6972 262868 6978 262880
rect 234246 262868 234252 262880
rect 6972 262840 234252 262868
rect 6972 262828 6978 262840
rect 234246 262828 234252 262840
rect 234304 262828 234310 262880
rect 234614 262828 234620 262880
rect 234672 262868 234678 262880
rect 283098 262868 283104 262880
rect 234672 262840 283104 262868
rect 234672 262828 234678 262840
rect 283098 262828 283104 262840
rect 283156 262828 283162 262880
rect 4798 259360 4804 259412
rect 4856 259400 4862 259412
rect 229094 259400 229100 259412
rect 4856 259372 229100 259400
rect 4856 259360 4862 259372
rect 229094 259360 229100 259372
rect 229152 259360 229158 259412
rect 354306 259360 354312 259412
rect 354364 259400 354370 259412
rect 580258 259400 580264 259412
rect 354364 259372 580264 259400
rect 354364 259360 354370 259372
rect 580258 259360 580264 259372
rect 580316 259360 580322 259412
rect 354122 258068 354128 258120
rect 354180 258108 354186 258120
rect 580166 258108 580172 258120
rect 354180 258080 580172 258108
rect 354180 258068 354186 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 229462 255252 229468 255264
rect 3476 255224 229468 255252
rect 3476 255212 3482 255224
rect 229462 255212 229468 255224
rect 229520 255212 229526 255264
rect 3510 251132 3516 251184
rect 3568 251172 3574 251184
rect 230382 251172 230388 251184
rect 3568 251144 230388 251172
rect 3568 251132 3574 251144
rect 230382 251132 230388 251144
rect 230440 251132 230446 251184
rect 353294 251132 353300 251184
rect 353352 251172 353358 251184
rect 360838 251172 360844 251184
rect 353352 251144 360844 251172
rect 353352 251132 353358 251144
rect 360838 251132 360844 251144
rect 360896 251132 360902 251184
rect 353294 248344 353300 248396
rect 353352 248384 353358 248396
rect 367738 248384 367744 248396
rect 353352 248356 367744 248384
rect 353352 248344 353358 248356
rect 367738 248344 367744 248356
rect 367796 248344 367802 248396
rect 32398 246984 32404 247036
rect 32456 247024 32462 247036
rect 229830 247024 229836 247036
rect 32456 246996 229836 247024
rect 32456 246984 32462 246996
rect 229830 246984 229836 246996
rect 229888 246984 229894 247036
rect 385678 244264 385684 244316
rect 385736 244304 385742 244316
rect 580166 244304 580172 244316
rect 385736 244276 580172 244304
rect 385736 244264 385742 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 353294 244196 353300 244248
rect 353352 244236 353358 244248
rect 374638 244236 374644 244248
rect 353352 244208 374644 244236
rect 353352 244196 353358 244208
rect 374638 244196 374644 244208
rect 374696 244196 374702 244248
rect 22738 242836 22744 242888
rect 22796 242876 22802 242888
rect 229646 242876 229652 242888
rect 22796 242848 229652 242876
rect 22796 242836 22802 242848
rect 229646 242836 229652 242848
rect 229704 242836 229710 242888
rect 353294 241408 353300 241460
rect 353352 241448 353358 241460
rect 381538 241448 381544 241460
rect 353352 241420 381544 241448
rect 353352 241408 353358 241420
rect 381538 241408 381544 241420
rect 381596 241408 381602 241460
rect 14458 240048 14464 240100
rect 14516 240088 14522 240100
rect 230382 240088 230388 240100
rect 14516 240060 230388 240088
rect 14516 240048 14522 240060
rect 230382 240048 230388 240060
rect 230440 240048 230446 240100
rect 353294 237328 353300 237380
rect 353352 237368 353358 237380
rect 580350 237368 580356 237380
rect 353352 237340 580356 237368
rect 353352 237328 353358 237340
rect 580350 237328 580356 237340
rect 580408 237328 580414 237380
rect 7558 235900 7564 235952
rect 7616 235940 7622 235952
rect 229830 235940 229836 235952
rect 7616 235912 229836 235940
rect 7616 235900 7622 235912
rect 229830 235900 229836 235912
rect 229888 235900 229894 235952
rect 353294 233180 353300 233232
rect 353352 233220 353358 233232
rect 580442 233220 580448 233232
rect 353352 233192 580448 233220
rect 353352 233180 353358 233192
rect 580442 233180 580448 233192
rect 580500 233180 580506 233232
rect 3602 231752 3608 231804
rect 3660 231792 3666 231804
rect 230382 231792 230388 231804
rect 3660 231764 230388 231792
rect 3660 231752 3666 231764
rect 230382 231752 230388 231764
rect 230440 231752 230446 231804
rect 353294 230392 353300 230444
rect 353352 230432 353358 230444
rect 359458 230432 359464 230444
rect 353352 230404 359464 230432
rect 353352 230392 353358 230404
rect 359458 230392 359464 230404
rect 359516 230392 359522 230444
rect 3694 227672 3700 227724
rect 3752 227712 3758 227724
rect 230382 227712 230388 227724
rect 3752 227684 230388 227712
rect 3752 227672 3758 227684
rect 230382 227672 230388 227684
rect 230440 227672 230446 227724
rect 353294 226244 353300 226296
rect 353352 226284 353358 226296
rect 364978 226284 364984 226296
rect 353352 226256 364984 226284
rect 353352 226244 353358 226256
rect 364978 226244 364984 226256
rect 365036 226244 365042 226296
rect 43438 224884 43444 224936
rect 43496 224924 43502 224936
rect 230382 224924 230388 224936
rect 43496 224896 230388 224924
rect 43496 224884 43502 224896
rect 230382 224884 230388 224896
rect 230440 224884 230446 224936
rect 353294 223524 353300 223576
rect 353352 223564 353358 223576
rect 373258 223564 373264 223576
rect 353352 223536 373264 223564
rect 353352 223524 353358 223536
rect 373258 223524 373264 223536
rect 373316 223524 373322 223576
rect 25498 220736 25504 220788
rect 25556 220776 25562 220788
rect 230382 220776 230388 220788
rect 25556 220748 230388 220776
rect 25556 220736 25562 220748
rect 230382 220736 230388 220748
rect 230440 220736 230446 220788
rect 353294 219308 353300 219360
rect 353352 219348 353358 219360
rect 356698 219348 356704 219360
rect 353352 219320 356704 219348
rect 353352 219308 353358 219320
rect 356698 219308 356704 219320
rect 356756 219308 356762 219360
rect 353938 218016 353944 218068
rect 353996 218056 354002 218068
rect 580166 218056 580172 218068
rect 353996 218028 580172 218056
rect 353996 218016 354002 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 17218 216588 17224 216640
rect 17276 216628 17282 216640
rect 230382 216628 230388 216640
rect 17276 216600 230388 216628
rect 17276 216588 17282 216600
rect 230382 216588 230388 216600
rect 230440 216588 230446 216640
rect 353294 216588 353300 216640
rect 353352 216628 353358 216640
rect 580442 216628 580448 216640
rect 353352 216600 580448 216628
rect 353352 216588 353358 216600
rect 580442 216588 580448 216600
rect 580500 216588 580506 216640
rect 8938 212440 8944 212492
rect 8996 212480 9002 212492
rect 230382 212480 230388 212492
rect 8996 212452 230388 212480
rect 8996 212440 9002 212452
rect 230382 212440 230388 212452
rect 230440 212440 230446 212492
rect 353294 212440 353300 212492
rect 353352 212480 353358 212492
rect 580626 212480 580632 212492
rect 353352 212452 580632 212480
rect 353352 212440 353358 212452
rect 580626 212440 580632 212452
rect 580684 212440 580690 212492
rect 3786 209720 3792 209772
rect 3844 209760 3850 209772
rect 230014 209760 230020 209772
rect 3844 209732 230020 209760
rect 3844 209720 3850 209732
rect 230014 209720 230020 209732
rect 230072 209720 230078 209772
rect 353294 209312 353300 209364
rect 353352 209352 353358 209364
rect 355318 209352 355324 209364
rect 353352 209324 355324 209352
rect 353352 209312 353358 209324
rect 355318 209312 355324 209324
rect 355376 209312 355382 209364
rect 3878 205572 3884 205624
rect 3936 205612 3942 205624
rect 230382 205612 230388 205624
rect 3936 205584 230388 205612
rect 3936 205572 3942 205584
rect 230382 205572 230388 205584
rect 230440 205572 230446 205624
rect 353294 205572 353300 205624
rect 353352 205612 353358 205624
rect 371878 205612 371884 205624
rect 353352 205584 371884 205612
rect 353352 205572 353358 205584
rect 371878 205572 371884 205584
rect 371936 205572 371942 205624
rect 31018 201424 31024 201476
rect 31076 201464 31082 201476
rect 229646 201464 229652 201476
rect 31076 201436 229652 201464
rect 31076 201424 31082 201436
rect 229646 201424 229652 201436
rect 229704 201424 229710 201476
rect 353294 201424 353300 201476
rect 353352 201464 353358 201476
rect 378778 201464 378784 201476
rect 353352 201436 378784 201464
rect 353352 201424 353358 201436
rect 378778 201424 378784 201436
rect 378836 201424 378842 201476
rect 353294 198636 353300 198688
rect 353352 198676 353358 198688
rect 363598 198676 363604 198688
rect 353352 198648 363604 198676
rect 353352 198636 353358 198648
rect 363598 198636 363604 198648
rect 363656 198636 363662 198688
rect 26878 197276 26884 197328
rect 26936 197316 26942 197328
rect 230382 197316 230388 197328
rect 26936 197288 230388 197316
rect 26936 197276 26942 197288
rect 230382 197276 230388 197288
rect 230440 197276 230446 197328
rect 18598 194488 18604 194540
rect 18656 194528 18662 194540
rect 229646 194528 229652 194540
rect 18656 194500 229652 194528
rect 18656 194488 18662 194500
rect 229646 194488 229652 194500
rect 229704 194488 229710 194540
rect 353294 194488 353300 194540
rect 353352 194528 353358 194540
rect 580718 194528 580724 194540
rect 353352 194500 580724 194528
rect 353352 194488 353358 194500
rect 580718 194488 580724 194500
rect 580776 194488 580782 194540
rect 10318 190408 10324 190460
rect 10376 190448 10382 190460
rect 230382 190448 230388 190460
rect 10376 190420 230388 190448
rect 10376 190408 10382 190420
rect 230382 190408 230388 190420
rect 230440 190408 230446 190460
rect 353294 187620 353300 187672
rect 353352 187660 353358 187672
rect 580810 187660 580816 187672
rect 353352 187632 580816 187660
rect 353352 187620 353358 187632
rect 580810 187620 580816 187632
rect 580868 187620 580874 187672
rect 3970 186260 3976 186312
rect 4028 186300 4034 186312
rect 230382 186300 230388 186312
rect 4028 186272 230388 186300
rect 4028 186260 4034 186272
rect 230382 186260 230388 186272
rect 230440 186260 230446 186312
rect 353294 183472 353300 183524
rect 353352 183512 353358 183524
rect 369118 183512 369124 183524
rect 353352 183484 369124 183512
rect 353352 183472 353358 183484
rect 369118 183472 369124 183484
rect 369176 183472 369182 183524
rect 4062 182112 4068 182164
rect 4120 182152 4126 182164
rect 230382 182152 230388 182164
rect 4120 182124 230388 182152
rect 4120 182112 4126 182124
rect 230382 182112 230388 182124
rect 230440 182112 230446 182164
rect 353294 180752 353300 180804
rect 353352 180792 353358 180804
rect 377398 180792 377404 180804
rect 353352 180764 377404 180792
rect 353352 180752 353358 180764
rect 377398 180752 377404 180764
rect 377456 180752 377462 180804
rect 221458 179324 221464 179376
rect 221516 179364 221522 179376
rect 229646 179364 229652 179376
rect 221516 179336 229652 179364
rect 221516 179324 221522 179336
rect 229646 179324 229652 179336
rect 229704 179324 229710 179376
rect 354030 178032 354036 178084
rect 354088 178072 354094 178084
rect 580166 178072 580172 178084
rect 354088 178044 580172 178072
rect 354088 178032 354094 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 353294 176604 353300 176656
rect 353352 176644 353358 176656
rect 442258 176644 442264 176656
rect 353352 176616 442264 176644
rect 353352 176604 353358 176616
rect 442258 176604 442264 176616
rect 442316 176604 442322 176656
rect 28258 175176 28264 175228
rect 28316 175216 28322 175228
rect 230382 175216 230388 175228
rect 28316 175188 230388 175216
rect 28316 175176 28322 175188
rect 230382 175176 230388 175188
rect 230440 175176 230446 175228
rect 353294 173816 353300 173868
rect 353352 173856 353358 173868
rect 580902 173856 580908 173868
rect 353352 173828 580908 173856
rect 353352 173816 353358 173828
rect 580902 173816 580908 173828
rect 580960 173816 580966 173868
rect 21358 171028 21364 171080
rect 21416 171068 21422 171080
rect 230382 171068 230388 171080
rect 21416 171040 230388 171068
rect 21416 171028 21422 171040
rect 230382 171028 230388 171040
rect 230440 171028 230446 171080
rect 13078 166948 13084 167000
rect 13136 166988 13142 167000
rect 230382 166988 230388 167000
rect 13136 166960 230388 166988
rect 13136 166948 13142 166960
rect 230382 166948 230388 166960
rect 230440 166948 230446 167000
rect 353294 166948 353300 167000
rect 353352 166988 353358 167000
rect 385678 166988 385684 167000
rect 353352 166960 385684 166988
rect 353352 166948 353358 166960
rect 385678 166948 385684 166960
rect 385736 166948 385742 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 229646 164200 229652 164212
rect 3384 164172 229652 164200
rect 3384 164160 3390 164172
rect 229646 164160 229652 164172
rect 229704 164160 229710 164212
rect 353294 162800 353300 162852
rect 353352 162840 353358 162852
rect 580258 162840 580264 162852
rect 353352 162812 580264 162840
rect 353352 162800 353358 162812
rect 580258 162800 580264 162812
rect 580316 162800 580322 162852
rect 3418 160012 3424 160064
rect 3476 160052 3482 160064
rect 229462 160052 229468 160064
rect 3476 160024 229468 160052
rect 3476 160012 3482 160024
rect 229462 160012 229468 160024
rect 229520 160012 229526 160064
rect 3510 155864 3516 155916
rect 3568 155904 3574 155916
rect 230382 155904 230388 155916
rect 3568 155876 230388 155904
rect 3568 155864 3574 155876
rect 230382 155864 230388 155876
rect 230440 155864 230446 155916
rect 353294 155864 353300 155916
rect 353352 155904 353358 155916
rect 580350 155904 580356 155916
rect 353352 155876 580356 155904
rect 353352 155864 353358 155876
rect 580350 155864 580356 155876
rect 580408 155864 580414 155916
rect 353938 151784 353944 151836
rect 353996 151824 354002 151836
rect 580166 151824 580172 151836
rect 353996 151796 580172 151824
rect 353996 151784 354002 151796
rect 580166 151784 580172 151796
rect 580224 151784 580230 151836
rect 3602 151716 3608 151768
rect 3660 151756 3666 151768
rect 230382 151756 230388 151768
rect 3660 151728 230388 151756
rect 3660 151716 3666 151728
rect 230382 151716 230388 151728
rect 230440 151716 230446 151768
rect 353294 151716 353300 151768
rect 353352 151756 353358 151768
rect 580442 151756 580448 151768
rect 353352 151728 580448 151756
rect 353352 151716 353358 151728
rect 580442 151716 580448 151728
rect 580500 151716 580506 151768
rect 3694 147568 3700 147620
rect 3752 147608 3758 147620
rect 229646 147608 229652 147620
rect 3752 147580 229652 147608
rect 3752 147568 3758 147580
rect 229646 147568 229652 147580
rect 229704 147568 229710 147620
rect 3786 144848 3792 144900
rect 3844 144888 3850 144900
rect 230382 144888 230388 144900
rect 3844 144860 230388 144888
rect 3844 144848 3850 144860
rect 230382 144848 230388 144860
rect 230440 144848 230446 144900
rect 353294 144848 353300 144900
rect 353352 144888 353358 144900
rect 580534 144888 580540 144900
rect 353352 144860 580540 144888
rect 353352 144848 353358 144860
rect 580534 144848 580540 144860
rect 580592 144848 580598 144900
rect 3418 140700 3424 140752
rect 3476 140740 3482 140752
rect 230382 140740 230388 140752
rect 3476 140712 230388 140740
rect 3476 140700 3482 140712
rect 230382 140700 230388 140712
rect 230440 140700 230446 140752
rect 353294 137980 353300 138032
rect 353352 138020 353358 138032
rect 580166 138020 580172 138032
rect 353352 137992 580172 138020
rect 353352 137980 353358 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 3418 136552 3424 136604
rect 3476 136592 3482 136604
rect 229830 136592 229836 136604
rect 3476 136564 229836 136592
rect 3476 136552 3482 136564
rect 229830 136552 229836 136564
rect 229888 136552 229894 136604
rect 3602 128324 3608 128376
rect 3660 128364 3666 128376
rect 230382 128364 230388 128376
rect 3660 128336 230388 128364
rect 3660 128324 3666 128336
rect 230382 128324 230388 128336
rect 230440 128324 230446 128376
rect 354306 126896 354312 126948
rect 354364 126936 354370 126948
rect 580166 126936 580172 126948
rect 354364 126908 580172 126936
rect 354364 126896 354370 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3510 115948 3516 116000
rect 3568 115988 3574 116000
rect 230198 115988 230204 116000
rect 3568 115960 230204 115988
rect 3568 115948 3574 115960
rect 230198 115948 230204 115960
rect 230256 115948 230262 116000
rect 353938 113092 353944 113144
rect 353996 113132 354002 113144
rect 579798 113132 579804 113144
rect 353996 113104 579804 113132
rect 353996 113092 354002 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 229738 111772 229744 111784
rect 3200 111744 229744 111772
rect 3200 111732 3206 111744
rect 229738 111732 229744 111744
rect 229796 111732 229802 111784
rect 3418 104864 3424 104916
rect 3476 104904 3482 104916
rect 230382 104904 230388 104916
rect 3476 104876 230388 104904
rect 3476 104864 3482 104876
rect 230382 104864 230388 104876
rect 230440 104864 230446 104916
rect 354582 100648 354588 100700
rect 354640 100688 354646 100700
rect 580166 100688 580172 100700
rect 354640 100660 580172 100688
rect 354640 100648 354646 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 238754 100104 238760 100156
rect 238812 100144 238818 100156
rect 239214 100144 239220 100156
rect 238812 100116 239220 100144
rect 238812 100104 238818 100116
rect 239214 100104 239220 100116
rect 239272 100104 239278 100156
rect 285674 100104 285680 100156
rect 285732 100144 285738 100156
rect 285950 100144 285956 100156
rect 285732 100116 285956 100144
rect 285732 100104 285738 100116
rect 285950 100104 285956 100116
rect 286008 100104 286014 100156
rect 225598 97928 225604 97980
rect 225656 97968 225662 97980
rect 276842 97968 276848 97980
rect 225656 97940 276848 97968
rect 225656 97928 225662 97940
rect 276842 97928 276848 97940
rect 276900 97928 276906 97980
rect 284938 97928 284944 97980
rect 284996 97968 285002 97980
rect 288802 97968 288808 97980
rect 284996 97940 288808 97968
rect 284996 97928 285002 97940
rect 288802 97928 288808 97940
rect 288860 97928 288866 97980
rect 334526 97928 334532 97980
rect 334584 97968 334590 97980
rect 336182 97968 336188 97980
rect 334584 97940 336188 97968
rect 334584 97928 334590 97940
rect 336182 97928 336188 97940
rect 336240 97928 336246 97980
rect 257154 97860 257160 97912
rect 257212 97900 257218 97912
rect 258626 97900 258632 97912
rect 257212 97872 258632 97900
rect 257212 97860 257218 97872
rect 258626 97860 258632 97872
rect 258684 97860 258690 97912
rect 268286 97792 268292 97844
rect 268344 97832 268350 97844
rect 281258 97832 281264 97844
rect 268344 97804 281264 97832
rect 268344 97792 268350 97804
rect 281258 97792 281264 97804
rect 281316 97792 281322 97844
rect 341794 97792 341800 97844
rect 341852 97832 341858 97844
rect 352558 97832 352564 97844
rect 341852 97804 352564 97832
rect 341852 97792 341858 97804
rect 352558 97792 352564 97804
rect 352616 97792 352622 97844
rect 224310 97724 224316 97776
rect 224368 97764 224374 97776
rect 241054 97764 241060 97776
rect 224368 97736 241060 97764
rect 224368 97724 224374 97736
rect 241054 97724 241060 97736
rect 241112 97724 241118 97776
rect 255958 97724 255964 97776
rect 256016 97764 256022 97776
rect 259362 97764 259368 97776
rect 256016 97736 259368 97764
rect 256016 97724 256022 97736
rect 259362 97724 259368 97736
rect 259420 97724 259426 97776
rect 275370 97724 275376 97776
rect 275428 97764 275434 97776
rect 279326 97764 279332 97776
rect 275428 97736 279332 97764
rect 275428 97724 275434 97736
rect 279326 97724 279332 97736
rect 279384 97724 279390 97776
rect 322106 97724 322112 97776
rect 322164 97764 322170 97776
rect 335630 97764 335636 97776
rect 322164 97736 335636 97764
rect 322164 97724 322170 97736
rect 335630 97724 335636 97736
rect 335688 97724 335694 97776
rect 349154 97724 349160 97776
rect 349212 97764 349218 97776
rect 364978 97764 364984 97776
rect 349212 97736 364984 97764
rect 349212 97724 349218 97736
rect 364978 97724 364984 97736
rect 365036 97724 365042 97776
rect 221458 97656 221464 97708
rect 221516 97696 221522 97708
rect 242526 97696 242532 97708
rect 221516 97668 242532 97696
rect 221516 97656 221522 97668
rect 242526 97656 242532 97668
rect 242584 97656 242590 97708
rect 345474 97656 345480 97708
rect 345532 97696 345538 97708
rect 363598 97696 363604 97708
rect 345532 97668 363604 97696
rect 345532 97656 345538 97668
rect 363598 97656 363604 97668
rect 363656 97656 363662 97708
rect 224218 97588 224224 97640
rect 224276 97628 224282 97640
rect 260282 97628 260288 97640
rect 224276 97600 260288 97628
rect 224276 97588 224282 97600
rect 260282 97588 260288 97600
rect 260340 97588 260346 97640
rect 266630 97628 266636 97640
rect 262324 97600 266636 97628
rect 228358 97520 228364 97572
rect 228416 97560 228422 97572
rect 262324 97560 262352 97600
rect 266630 97588 266636 97600
rect 266688 97588 266694 97640
rect 274358 97588 274364 97640
rect 274416 97628 274422 97640
rect 281718 97628 281724 97640
rect 274416 97600 281724 97628
rect 274416 97588 274422 97600
rect 281718 97588 281724 97600
rect 281776 97588 281782 97640
rect 294414 97588 294420 97640
rect 294472 97628 294478 97640
rect 302234 97628 302240 97640
rect 294472 97600 302240 97628
rect 294472 97588 294478 97600
rect 302234 97588 302240 97600
rect 302292 97588 302298 97640
rect 317046 97588 317052 97640
rect 317104 97628 317110 97640
rect 333330 97628 333336 97640
rect 317104 97600 333336 97628
rect 317104 97588 317110 97600
rect 333330 97588 333336 97600
rect 333388 97588 333394 97640
rect 335906 97588 335912 97640
rect 335964 97628 335970 97640
rect 355318 97628 355324 97640
rect 335964 97600 355324 97628
rect 335964 97588 335970 97600
rect 355318 97588 355324 97600
rect 355376 97588 355382 97640
rect 228416 97532 262352 97560
rect 228416 97520 228422 97532
rect 275278 97520 275284 97572
rect 275336 97560 275342 97572
rect 283466 97560 283472 97572
rect 275336 97532 283472 97560
rect 275336 97520 275342 97532
rect 283466 97520 283472 97532
rect 283524 97520 283530 97572
rect 295610 97520 295616 97572
rect 295668 97560 295674 97572
rect 307202 97560 307208 97572
rect 295668 97532 307208 97560
rect 295668 97520 295674 97532
rect 307202 97520 307208 97532
rect 307260 97520 307266 97572
rect 311894 97520 311900 97572
rect 311952 97560 311958 97572
rect 332134 97560 332140 97572
rect 311952 97532 332140 97560
rect 311952 97520 311958 97532
rect 332134 97520 332140 97532
rect 332192 97520 332198 97572
rect 338206 97520 338212 97572
rect 338264 97560 338270 97572
rect 360838 97560 360844 97572
rect 338264 97532 360844 97560
rect 338264 97520 338270 97532
rect 360838 97520 360844 97532
rect 360896 97520 360902 97572
rect 295334 97452 295340 97504
rect 295392 97492 295398 97504
rect 307018 97492 307024 97504
rect 295392 97464 307024 97492
rect 295392 97452 295398 97464
rect 307018 97452 307024 97464
rect 307076 97452 307082 97504
rect 330846 97452 330852 97504
rect 330904 97492 330910 97504
rect 355502 97492 355508 97504
rect 330904 97464 355508 97492
rect 330904 97452 330910 97464
rect 355502 97452 355508 97464
rect 355560 97452 355566 97504
rect 124214 97384 124220 97436
rect 124272 97424 124278 97436
rect 257614 97424 257620 97436
rect 124272 97396 257620 97424
rect 124272 97384 124278 97396
rect 257614 97384 257620 97396
rect 257672 97384 257678 97436
rect 276658 97384 276664 97436
rect 276716 97424 276722 97436
rect 278038 97424 278044 97436
rect 276716 97396 278044 97424
rect 276716 97384 276722 97396
rect 278038 97384 278044 97396
rect 278096 97384 278102 97436
rect 279418 97384 279424 97436
rect 279476 97424 279482 97436
rect 288526 97424 288532 97436
rect 279476 97396 288532 97424
rect 279476 97384 279482 97396
rect 288526 97384 288532 97396
rect 288584 97384 288590 97436
rect 297266 97384 297272 97436
rect 297324 97424 297330 97436
rect 311158 97424 311164 97436
rect 297324 97396 311164 97424
rect 297324 97384 297330 97396
rect 311158 97384 311164 97396
rect 311216 97384 311222 97436
rect 331582 97384 331588 97436
rect 331640 97424 331646 97436
rect 356698 97424 356704 97436
rect 331640 97396 356704 97424
rect 331640 97384 331646 97396
rect 356698 97384 356704 97396
rect 356756 97384 356762 97436
rect 106274 97316 106280 97368
rect 106332 97356 106338 97368
rect 254026 97356 254032 97368
rect 106332 97328 254032 97356
rect 106332 97316 106338 97328
rect 254026 97316 254032 97328
rect 254084 97316 254090 97368
rect 269758 97316 269764 97368
rect 269816 97356 269822 97368
rect 280798 97356 280804 97368
rect 269816 97328 280804 97356
rect 269816 97316 269822 97328
rect 280798 97316 280804 97328
rect 280856 97316 280862 97368
rect 300946 97316 300952 97368
rect 301004 97356 301010 97368
rect 331858 97356 331864 97368
rect 301004 97328 331864 97356
rect 301004 97316 301010 97328
rect 331858 97316 331864 97328
rect 331916 97316 331922 97368
rect 335262 97316 335268 97368
rect 335320 97356 335326 97368
rect 359458 97356 359464 97368
rect 335320 97328 359464 97356
rect 335320 97316 335326 97328
rect 359458 97316 359464 97328
rect 359516 97316 359522 97368
rect 10318 97248 10324 97300
rect 10376 97288 10382 97300
rect 233050 97288 233056 97300
rect 10376 97260 233056 97288
rect 10376 97248 10382 97260
rect 233050 97248 233056 97260
rect 233108 97248 233114 97300
rect 257338 97248 257344 97300
rect 257396 97288 257402 97300
rect 265158 97288 265164 97300
rect 257396 97260 265164 97288
rect 257396 97248 257402 97260
rect 265158 97248 265164 97260
rect 265216 97248 265222 97300
rect 298738 97248 298744 97300
rect 298796 97288 298802 97300
rect 319438 97288 319444 97300
rect 298796 97260 319444 97288
rect 298796 97248 298802 97260
rect 319438 97248 319444 97260
rect 319496 97248 319502 97300
rect 332318 97248 332324 97300
rect 332376 97288 332382 97300
rect 485038 97288 485044 97300
rect 332376 97260 485044 97288
rect 332376 97248 332382 97260
rect 485038 97248 485044 97260
rect 485096 97248 485102 97300
rect 303706 97180 303712 97232
rect 303764 97220 303770 97232
rect 304442 97220 304448 97232
rect 303764 97192 304448 97220
rect 303764 97180 303770 97192
rect 304442 97180 304448 97192
rect 304500 97180 304506 97232
rect 350810 97112 350816 97164
rect 350868 97152 350874 97164
rect 355410 97152 355416 97164
rect 350868 97124 355416 97152
rect 350868 97112 350874 97124
rect 355410 97112 355416 97124
rect 355468 97112 355474 97164
rect 242986 97044 242992 97096
rect 243044 97084 243050 97096
rect 244734 97084 244740 97096
rect 243044 97056 244740 97084
rect 243044 97044 243050 97056
rect 244734 97044 244740 97056
rect 244792 97044 244798 97096
rect 279142 97044 279148 97096
rect 279200 97084 279206 97096
rect 279878 97084 279884 97096
rect 279200 97056 279884 97084
rect 279200 97044 279206 97056
rect 279878 97044 279884 97056
rect 279936 97044 279942 97096
rect 295426 97044 295432 97096
rect 295484 97084 295490 97096
rect 295886 97084 295892 97096
rect 295484 97056 295892 97084
rect 295484 97044 295490 97056
rect 295886 97044 295892 97056
rect 295944 97044 295950 97096
rect 296898 97044 296904 97096
rect 296956 97084 296962 97096
rect 297358 97084 297364 97096
rect 296956 97056 297364 97084
rect 296956 97044 296962 97056
rect 297358 97044 297364 97056
rect 297416 97044 297422 97096
rect 301038 97044 301044 97096
rect 301096 97084 301102 97096
rect 301498 97084 301504 97096
rect 301096 97056 301504 97084
rect 301096 97044 301102 97056
rect 301498 97044 301504 97056
rect 301556 97044 301562 97096
rect 303706 97044 303712 97096
rect 303764 97084 303770 97096
rect 304166 97084 304172 97096
rect 303764 97056 304172 97084
rect 303764 97044 303770 97056
rect 304166 97044 304172 97056
rect 304224 97044 304230 97096
rect 305178 97044 305184 97096
rect 305236 97084 305242 97096
rect 305638 97084 305644 97096
rect 305236 97056 305644 97084
rect 305236 97044 305242 97056
rect 305638 97044 305644 97056
rect 305696 97044 305702 97096
rect 327074 97044 327080 97096
rect 327132 97084 327138 97096
rect 327534 97084 327540 97096
rect 327132 97056 327540 97084
rect 327132 97044 327138 97056
rect 327534 97044 327540 97056
rect 327592 97044 327598 97096
rect 328546 97044 328552 97096
rect 328604 97084 328610 97096
rect 329006 97084 329012 97096
rect 328604 97056 329012 97084
rect 328604 97044 328610 97056
rect 329006 97044 329012 97056
rect 329064 97044 329070 97096
rect 231118 96976 231124 97028
rect 231176 97016 231182 97028
rect 233510 97016 233516 97028
rect 231176 96988 233516 97016
rect 231176 96976 231182 96988
rect 233510 96976 233516 96988
rect 233568 96976 233574 97028
rect 233878 96976 233884 97028
rect 233936 97016 233942 97028
rect 236454 97016 236460 97028
rect 233936 96988 236460 97016
rect 233936 96976 233942 96988
rect 236454 96976 236460 96988
rect 236512 96976 236518 97028
rect 278038 96976 278044 97028
rect 278096 97016 278102 97028
rect 280522 97016 280528 97028
rect 278096 96988 280528 97016
rect 278096 96976 278102 96988
rect 280522 96976 280528 96988
rect 280580 96976 280586 97028
rect 298278 96976 298284 97028
rect 298336 97016 298342 97028
rect 305730 97016 305736 97028
rect 298336 96988 305736 97016
rect 298336 96976 298342 96988
rect 305730 96976 305736 96988
rect 305788 96976 305794 97028
rect 325786 96976 325792 97028
rect 325844 97016 325850 97028
rect 327718 97016 327724 97028
rect 325844 96988 327724 97016
rect 325844 96976 325850 96988
rect 327718 96976 327724 96988
rect 327776 96976 327782 97028
rect 328730 96976 328736 97028
rect 328788 97016 328794 97028
rect 333238 97016 333244 97028
rect 328788 96988 333244 97016
rect 328788 96976 328794 96988
rect 333238 96976 333244 96988
rect 333296 96976 333302 97028
rect 348418 96976 348424 97028
rect 348476 97016 348482 97028
rect 352742 97016 352748 97028
rect 348476 96988 352748 97016
rect 348476 96976 348482 96988
rect 352742 96976 352748 96988
rect 352800 96976 352806 97028
rect 231946 96908 231952 96960
rect 232004 96948 232010 96960
rect 232774 96948 232780 96960
rect 232004 96920 232780 96948
rect 232004 96908 232010 96920
rect 232774 96908 232780 96920
rect 232832 96908 232838 96960
rect 233602 96908 233608 96960
rect 233660 96948 233666 96960
rect 234246 96948 234252 96960
rect 233660 96920 234252 96948
rect 233660 96908 233666 96920
rect 234246 96908 234252 96920
rect 234304 96908 234310 96960
rect 234614 96908 234620 96960
rect 234672 96948 234678 96960
rect 235350 96948 235356 96960
rect 234672 96920 235356 96948
rect 234672 96908 234678 96920
rect 235350 96908 235356 96920
rect 235408 96908 235414 96960
rect 237742 96908 237748 96960
rect 237800 96948 237806 96960
rect 238018 96948 238024 96960
rect 237800 96920 238024 96948
rect 237800 96908 237806 96920
rect 238018 96908 238024 96920
rect 238076 96908 238082 96960
rect 239398 96908 239404 96960
rect 239456 96948 239462 96960
rect 240318 96948 240324 96960
rect 239456 96920 240324 96948
rect 239456 96908 239462 96920
rect 240318 96908 240324 96920
rect 240376 96908 240382 96960
rect 242158 96908 242164 96960
rect 242216 96948 242222 96960
rect 245470 96948 245476 96960
rect 242216 96920 245476 96948
rect 242216 96908 242222 96920
rect 245470 96908 245476 96920
rect 245528 96908 245534 96960
rect 255774 96908 255780 96960
rect 255832 96948 255838 96960
rect 256142 96948 256148 96960
rect 255832 96920 256148 96948
rect 255832 96908 255838 96920
rect 256142 96908 256148 96920
rect 256200 96908 256206 96960
rect 256970 96908 256976 96960
rect 257028 96948 257034 96960
rect 257246 96948 257252 96960
rect 257028 96920 257252 96948
rect 257028 96908 257034 96920
rect 257246 96908 257252 96920
rect 257304 96908 257310 96960
rect 259914 96908 259920 96960
rect 259972 96948 259978 96960
rect 260374 96948 260380 96960
rect 259972 96920 260380 96948
rect 259972 96908 259978 96920
rect 260374 96908 260380 96920
rect 260432 96908 260438 96960
rect 261110 96908 261116 96960
rect 261168 96948 261174 96960
rect 261386 96948 261392 96960
rect 261168 96920 261392 96948
rect 261168 96908 261174 96920
rect 261386 96908 261392 96920
rect 261444 96908 261450 96960
rect 262582 96908 262588 96960
rect 262640 96948 262646 96960
rect 263318 96948 263324 96960
rect 262640 96920 263324 96948
rect 262640 96908 262646 96920
rect 263318 96908 263324 96920
rect 263376 96908 263382 96960
rect 275462 96908 275468 96960
rect 275520 96948 275526 96960
rect 276106 96948 276112 96960
rect 275520 96920 276112 96948
rect 275520 96908 275526 96920
rect 276106 96908 276112 96920
rect 276164 96908 276170 96960
rect 276198 96908 276204 96960
rect 276256 96948 276262 96960
rect 277302 96948 277308 96960
rect 276256 96920 277308 96948
rect 276256 96908 276262 96920
rect 277302 96908 277308 96920
rect 277360 96908 277366 96960
rect 279602 96908 279608 96960
rect 279660 96948 279666 96960
rect 279878 96948 279884 96960
rect 279660 96920 279884 96948
rect 279660 96908 279666 96920
rect 279878 96908 279884 96920
rect 279936 96908 279942 96960
rect 281810 96908 281816 96960
rect 281868 96948 281874 96960
rect 282178 96948 282184 96960
rect 281868 96920 282184 96948
rect 281868 96908 281874 96920
rect 282178 96908 282184 96920
rect 282236 96908 282242 96960
rect 283282 96908 283288 96960
rect 283340 96948 283346 96960
rect 284018 96948 284024 96960
rect 283340 96920 284024 96948
rect 283340 96908 283346 96920
rect 284018 96908 284024 96920
rect 284076 96908 284082 96960
rect 284662 96908 284668 96960
rect 284720 96948 284726 96960
rect 285214 96948 285220 96960
rect 284720 96920 285220 96948
rect 284720 96908 284726 96920
rect 285214 96908 285220 96920
rect 285272 96908 285278 96960
rect 286410 96908 286416 96960
rect 286468 96948 286474 96960
rect 286686 96948 286692 96960
rect 286468 96920 286692 96948
rect 286468 96908 286474 96920
rect 286686 96908 286692 96920
rect 286744 96908 286750 96960
rect 287146 96908 287152 96960
rect 287204 96948 287210 96960
rect 287422 96948 287428 96960
rect 287204 96920 287428 96948
rect 287204 96908 287210 96920
rect 287422 96908 287428 96920
rect 287480 96908 287486 96960
rect 287882 96908 287888 96960
rect 287940 96948 287946 96960
rect 288158 96948 288164 96960
rect 287940 96920 288164 96948
rect 287940 96908 287946 96920
rect 288158 96908 288164 96920
rect 288216 96908 288222 96960
rect 290090 96908 290096 96960
rect 290148 96948 290154 96960
rect 290826 96948 290832 96960
rect 290148 96920 290832 96948
rect 290148 96908 290154 96920
rect 290826 96908 290832 96920
rect 290884 96908 290890 96960
rect 291562 96908 291568 96960
rect 291620 96948 291626 96960
rect 292390 96948 292396 96960
rect 291620 96920 292396 96948
rect 291620 96908 291626 96920
rect 292390 96908 292396 96920
rect 292448 96908 292454 96960
rect 292758 96908 292764 96960
rect 292816 96948 292822 96960
rect 293126 96948 293132 96960
rect 292816 96920 293132 96948
rect 292816 96908 292822 96920
rect 293126 96908 293132 96920
rect 293184 96908 293190 96960
rect 294230 96908 294236 96960
rect 294288 96948 294294 96960
rect 294690 96948 294696 96960
rect 294288 96920 294696 96948
rect 294288 96908 294294 96920
rect 294690 96908 294696 96920
rect 294748 96908 294754 96960
rect 295886 96908 295892 96960
rect 295944 96948 295950 96960
rect 296530 96948 296536 96960
rect 295944 96920 296536 96948
rect 295944 96908 295950 96920
rect 296530 96908 296536 96920
rect 296588 96908 296594 96960
rect 297358 96908 297364 96960
rect 297416 96948 297422 96960
rect 298002 96948 298008 96960
rect 297416 96920 298008 96948
rect 297416 96908 297422 96920
rect 298002 96908 298008 96920
rect 298060 96908 298066 96960
rect 298370 96908 298376 96960
rect 298428 96948 298434 96960
rect 298830 96948 298836 96960
rect 298428 96920 298836 96948
rect 298428 96908 298434 96920
rect 298830 96908 298836 96920
rect 298888 96908 298894 96960
rect 299566 96908 299572 96960
rect 299624 96948 299630 96960
rect 299934 96948 299940 96960
rect 299624 96920 299940 96948
rect 299624 96908 299630 96920
rect 299934 96908 299940 96920
rect 299992 96908 299998 96960
rect 300026 96908 300032 96960
rect 300084 96948 300090 96960
rect 300670 96948 300676 96960
rect 300084 96920 300676 96948
rect 300084 96908 300090 96920
rect 300670 96908 300676 96920
rect 300728 96908 300734 96960
rect 302510 96908 302516 96960
rect 302568 96948 302574 96960
rect 302970 96948 302976 96960
rect 302568 96920 302976 96948
rect 302568 96908 302574 96920
rect 302970 96908 302976 96920
rect 303028 96908 303034 96960
rect 304166 96908 304172 96960
rect 304224 96948 304230 96960
rect 304810 96948 304816 96960
rect 304224 96920 304816 96948
rect 304224 96908 304230 96920
rect 304810 96908 304816 96920
rect 304868 96908 304874 96960
rect 305638 96908 305644 96960
rect 305696 96948 305702 96960
rect 306282 96948 306288 96960
rect 305696 96920 306288 96948
rect 305696 96908 305702 96920
rect 306282 96908 306288 96920
rect 306340 96908 306346 96960
rect 306650 96908 306656 96960
rect 306708 96948 306714 96960
rect 307478 96948 307484 96960
rect 306708 96920 307484 96948
rect 306708 96908 306714 96920
rect 307478 96908 307484 96920
rect 307536 96908 307542 96960
rect 307846 96908 307852 96960
rect 307904 96948 307910 96960
rect 308582 96948 308588 96960
rect 307904 96920 308588 96948
rect 307904 96908 307910 96920
rect 308582 96908 308588 96920
rect 308640 96908 308646 96960
rect 309318 96908 309324 96960
rect 309376 96948 309382 96960
rect 310054 96948 310060 96960
rect 309376 96920 310060 96948
rect 309376 96908 309382 96920
rect 310054 96908 310060 96920
rect 310112 96908 310118 96960
rect 310514 96908 310520 96960
rect 310572 96948 310578 96960
rect 310882 96948 310888 96960
rect 310572 96920 310888 96948
rect 310572 96908 310578 96920
rect 310882 96908 310888 96920
rect 310940 96908 310946 96960
rect 312446 96908 312452 96960
rect 312504 96948 312510 96960
rect 312722 96948 312728 96960
rect 312504 96920 312728 96948
rect 312504 96908 312510 96920
rect 312722 96908 312728 96920
rect 312780 96908 312786 96960
rect 313458 96908 313464 96960
rect 313516 96948 313522 96960
rect 313826 96948 313832 96960
rect 313516 96920 313832 96948
rect 313516 96908 313522 96920
rect 313826 96908 313832 96920
rect 313884 96908 313890 96960
rect 313918 96908 313924 96960
rect 313976 96948 313982 96960
rect 314194 96948 314200 96960
rect 313976 96920 314200 96948
rect 313976 96908 313982 96920
rect 314194 96908 314200 96920
rect 314252 96908 314258 96960
rect 314654 96908 314660 96960
rect 314712 96948 314718 96960
rect 315758 96948 315764 96960
rect 314712 96920 315764 96948
rect 314712 96908 314718 96920
rect 315758 96908 315764 96920
rect 315816 96908 315822 96960
rect 316126 96908 316132 96960
rect 316184 96948 316190 96960
rect 316586 96948 316592 96960
rect 316184 96920 316592 96948
rect 316184 96908 316190 96920
rect 316586 96908 316592 96920
rect 316644 96908 316650 96960
rect 317598 96908 317604 96960
rect 317656 96948 317662 96960
rect 318518 96948 318524 96960
rect 317656 96920 318524 96948
rect 317656 96908 317662 96920
rect 318518 96908 318524 96920
rect 318576 96908 318582 96960
rect 318794 96908 318800 96960
rect 318852 96948 318858 96960
rect 319530 96948 319536 96960
rect 318852 96920 319536 96948
rect 318852 96908 318858 96920
rect 319530 96908 319536 96920
rect 319588 96908 319594 96960
rect 321738 96908 321744 96960
rect 321796 96948 321802 96960
rect 322566 96948 322572 96960
rect 321796 96920 322572 96948
rect 321796 96908 321802 96920
rect 322566 96908 322572 96920
rect 322624 96908 322630 96960
rect 322934 96908 322940 96960
rect 322992 96948 322998 96960
rect 323302 96948 323308 96960
rect 322992 96920 323308 96948
rect 322992 96908 322998 96920
rect 323302 96908 323308 96920
rect 323360 96908 323366 96960
rect 323394 96908 323400 96960
rect 323452 96948 323458 96960
rect 324038 96948 324044 96960
rect 323452 96920 324044 96948
rect 323452 96908 323458 96920
rect 324038 96908 324044 96920
rect 324096 96908 324102 96960
rect 324406 96908 324412 96960
rect 324464 96948 324470 96960
rect 325510 96948 325516 96960
rect 324464 96920 325516 96948
rect 324464 96908 324470 96920
rect 325510 96908 325516 96920
rect 325568 96908 325574 96960
rect 327534 96908 327540 96960
rect 327592 96948 327598 96960
rect 328178 96948 328184 96960
rect 327592 96920 328184 96948
rect 327592 96908 327598 96920
rect 328178 96908 328184 96920
rect 328236 96908 328242 96960
rect 329006 96908 329012 96960
rect 329064 96948 329070 96960
rect 329650 96948 329656 96960
rect 329064 96920 329656 96948
rect 329064 96908 329070 96920
rect 329650 96908 329656 96920
rect 329708 96908 329714 96960
rect 330202 96908 330208 96960
rect 330260 96948 330266 96960
rect 330478 96948 330484 96960
rect 330260 96920 330484 96948
rect 330260 96908 330266 96920
rect 330478 96908 330484 96920
rect 330536 96908 330542 96960
rect 332686 96908 332692 96960
rect 332744 96948 332750 96960
rect 333514 96948 333520 96960
rect 332744 96920 333520 96948
rect 332744 96908 332750 96920
rect 333514 96908 333520 96920
rect 333572 96908 333578 96960
rect 334342 96908 334348 96960
rect 334400 96948 334406 96960
rect 334986 96948 334992 96960
rect 334400 96920 334992 96948
rect 334400 96908 334406 96920
rect 334986 96908 334992 96920
rect 335044 96908 335050 96960
rect 335354 96908 335360 96960
rect 335412 96948 335418 96960
rect 336458 96948 336464 96960
rect 335412 96920 336464 96948
rect 335412 96908 335418 96920
rect 336458 96908 336464 96920
rect 336516 96908 336522 96960
rect 337286 96908 337292 96960
rect 337344 96948 337350 96960
rect 337654 96948 337660 96960
rect 337344 96920 337660 96948
rect 337344 96908 337350 96920
rect 337654 96908 337660 96920
rect 337712 96908 337718 96960
rect 338758 96908 338764 96960
rect 338816 96948 338822 96960
rect 339218 96948 339224 96960
rect 338816 96920 339224 96948
rect 338816 96908 338822 96920
rect 339218 96908 339224 96920
rect 339276 96908 339282 96960
rect 339494 96908 339500 96960
rect 339552 96948 339558 96960
rect 339862 96948 339868 96960
rect 339552 96920 339868 96948
rect 339552 96908 339558 96920
rect 339862 96908 339868 96920
rect 339920 96908 339926 96960
rect 339954 96908 339960 96960
rect 340012 96948 340018 96960
rect 340598 96948 340604 96960
rect 340012 96920 340604 96948
rect 340012 96908 340018 96920
rect 340598 96908 340604 96920
rect 340656 96908 340662 96960
rect 341150 96908 341156 96960
rect 341208 96948 341214 96960
rect 341426 96948 341432 96960
rect 341208 96920 341432 96948
rect 341208 96908 341214 96920
rect 341426 96908 341432 96920
rect 341484 96908 341490 96960
rect 342622 96908 342628 96960
rect 342680 96948 342686 96960
rect 343358 96948 343364 96960
rect 342680 96920 343364 96948
rect 342680 96908 342686 96920
rect 343358 96908 343364 96920
rect 343416 96908 343422 96960
rect 344094 96908 344100 96960
rect 344152 96948 344158 96960
rect 344738 96948 344744 96960
rect 344152 96920 344744 96948
rect 344152 96908 344158 96920
rect 344738 96908 344744 96920
rect 344796 96908 344802 96960
rect 345290 96908 345296 96960
rect 345348 96948 345354 96960
rect 345934 96948 345940 96960
rect 345348 96920 345940 96948
rect 345348 96908 345354 96920
rect 345934 96908 345940 96920
rect 345992 96908 345998 96960
rect 346762 96908 346768 96960
rect 346820 96948 346826 96960
rect 347406 96948 347412 96960
rect 346820 96920 347412 96948
rect 346820 96908 346826 96920
rect 347406 96908 347412 96920
rect 347464 96908 347470 96960
rect 347774 96908 347780 96960
rect 347832 96948 347838 96960
rect 348602 96948 348608 96960
rect 347832 96920 348608 96948
rect 347832 96908 347838 96920
rect 348602 96908 348608 96920
rect 348660 96908 348666 96960
rect 349706 96908 349712 96960
rect 349764 96948 349770 96960
rect 350166 96948 350172 96960
rect 349764 96920 350172 96948
rect 349764 96908 349770 96920
rect 350166 96908 350172 96920
rect 350224 96908 350230 96960
rect 350902 96908 350908 96960
rect 350960 96948 350966 96960
rect 351178 96948 351184 96960
rect 350960 96920 351184 96948
rect 350960 96908 350966 96920
rect 351178 96908 351184 96920
rect 351236 96908 351242 96960
rect 235258 96840 235264 96892
rect 235316 96880 235322 96892
rect 236730 96880 236736 96892
rect 235316 96852 236736 96880
rect 235316 96840 235322 96852
rect 236730 96840 236736 96852
rect 236788 96840 236794 96892
rect 240134 96840 240140 96892
rect 240192 96880 240198 96892
rect 241422 96880 241428 96892
rect 240192 96852 241428 96880
rect 240192 96840 240198 96852
rect 241422 96840 241428 96852
rect 241480 96840 241486 96892
rect 243354 96840 243360 96892
rect 243412 96880 243418 96892
rect 243722 96880 243728 96892
rect 243412 96852 243728 96880
rect 243412 96840 243418 96852
rect 243722 96840 243728 96852
rect 243780 96840 243786 96892
rect 255498 96840 255504 96892
rect 255556 96880 255562 96892
rect 256234 96880 256240 96892
rect 255556 96852 256240 96880
rect 255556 96840 255562 96852
rect 256234 96840 256240 96852
rect 256292 96840 256298 96892
rect 260098 96840 260104 96892
rect 260156 96880 260162 96892
rect 261018 96880 261024 96892
rect 260156 96852 261024 96880
rect 260156 96840 260162 96852
rect 261018 96840 261024 96852
rect 261076 96840 261082 96892
rect 261478 96840 261484 96892
rect 261536 96880 261542 96892
rect 262950 96880 262956 96892
rect 261536 96852 262956 96880
rect 261536 96840 261542 96852
rect 262950 96840 262956 96852
rect 263008 96840 263014 96892
rect 270494 96840 270500 96892
rect 270552 96880 270558 96892
rect 272518 96880 272524 96892
rect 270552 96852 272524 96880
rect 270552 96840 270558 96852
rect 272518 96840 272524 96852
rect 272576 96840 272582 96892
rect 275002 96840 275008 96892
rect 275060 96880 275066 96892
rect 275738 96880 275744 96892
rect 275060 96852 275744 96880
rect 275060 96840 275066 96852
rect 275738 96840 275744 96852
rect 275796 96840 275802 96892
rect 279510 96840 279516 96892
rect 279568 96880 279574 96892
rect 280246 96880 280252 96892
rect 279568 96852 280252 96880
rect 279568 96840 279574 96852
rect 280246 96840 280252 96852
rect 280304 96840 280310 96892
rect 287238 96840 287244 96892
rect 287296 96840 287302 96892
rect 289078 96840 289084 96892
rect 289136 96880 289142 96892
rect 289998 96880 290004 96892
rect 289136 96852 290004 96880
rect 289136 96840 289142 96852
rect 289998 96840 290004 96852
rect 290056 96840 290062 96892
rect 298094 96840 298100 96892
rect 298152 96880 298158 96892
rect 299106 96880 299112 96892
rect 298152 96852 299112 96880
rect 298152 96840 298158 96852
rect 299106 96840 299112 96852
rect 299164 96840 299170 96892
rect 306374 96840 306380 96892
rect 306432 96880 306438 96892
rect 307110 96880 307116 96892
rect 306432 96852 307116 96880
rect 306432 96840 306438 96852
rect 307110 96840 307116 96852
rect 307168 96840 307174 96892
rect 311986 96840 311992 96892
rect 312044 96880 312050 96892
rect 313090 96880 313096 96892
rect 312044 96852 313096 96880
rect 312044 96840 312050 96852
rect 313090 96840 313096 96852
rect 313148 96840 313154 96892
rect 336826 96840 336832 96892
rect 336884 96880 336890 96892
rect 337746 96880 337752 96892
rect 336884 96852 337752 96880
rect 336884 96840 336890 96852
rect 337746 96840 337752 96852
rect 337804 96840 337810 96892
rect 338482 96840 338488 96892
rect 338540 96880 338546 96892
rect 339126 96880 339132 96892
rect 338540 96852 339132 96880
rect 338540 96840 338546 96852
rect 339126 96840 339132 96852
rect 339184 96840 339190 96892
rect 343634 96840 343640 96892
rect 343692 96880 343698 96892
rect 344370 96880 344376 96892
rect 343692 96852 344376 96880
rect 343692 96840 343698 96852
rect 344370 96840 344376 96852
rect 344428 96840 344434 96892
rect 349430 96840 349436 96892
rect 349488 96880 349494 96892
rect 350074 96880 350080 96892
rect 349488 96852 350080 96880
rect 349488 96840 349494 96852
rect 350074 96840 350080 96852
rect 350132 96840 350138 96892
rect 350626 96840 350632 96892
rect 350684 96880 350690 96892
rect 352650 96880 352656 96892
rect 350684 96852 352656 96880
rect 350684 96840 350690 96852
rect 352650 96840 352656 96852
rect 352708 96840 352714 96892
rect 238018 96772 238024 96824
rect 238076 96812 238082 96824
rect 238478 96812 238484 96824
rect 238076 96784 238484 96812
rect 238076 96772 238082 96784
rect 238478 96772 238484 96784
rect 238536 96772 238542 96824
rect 243538 96772 243544 96824
rect 243596 96812 243602 96824
rect 244274 96812 244280 96824
rect 243596 96784 244280 96812
rect 243596 96772 243602 96784
rect 244274 96772 244280 96784
rect 244332 96772 244338 96824
rect 261386 96772 261392 96824
rect 261444 96812 261450 96824
rect 261846 96812 261852 96824
rect 261444 96784 261852 96812
rect 261444 96772 261450 96784
rect 261846 96772 261852 96784
rect 261904 96772 261910 96824
rect 273990 96772 273996 96824
rect 274048 96812 274054 96824
rect 274910 96812 274916 96824
rect 274048 96784 274916 96812
rect 274048 96772 274054 96784
rect 274910 96772 274916 96784
rect 274968 96772 274974 96824
rect 280798 96772 280804 96824
rect 280856 96812 280862 96824
rect 284386 96812 284392 96824
rect 280856 96784 284392 96812
rect 280856 96772 280862 96784
rect 284386 96772 284392 96784
rect 284444 96772 284450 96824
rect 232498 96704 232504 96756
rect 232556 96744 232562 96756
rect 234522 96744 234528 96756
rect 232556 96716 234528 96744
rect 232556 96704 232562 96716
rect 234522 96704 234528 96716
rect 234580 96704 234586 96756
rect 260190 96704 260196 96756
rect 260248 96744 260254 96756
rect 262214 96744 262220 96756
rect 260248 96716 262220 96744
rect 260248 96704 260254 96716
rect 262214 96704 262220 96716
rect 262272 96704 262278 96756
rect 265434 96704 265440 96756
rect 265492 96744 265498 96756
rect 267366 96744 267372 96756
rect 265492 96716 267372 96744
rect 265492 96704 265498 96716
rect 267366 96704 267372 96716
rect 267424 96704 267430 96756
rect 282178 96704 282184 96756
rect 282236 96744 282242 96756
rect 283190 96744 283196 96756
rect 282236 96716 283196 96744
rect 282236 96704 282242 96716
rect 283190 96704 283196 96716
rect 283248 96704 283254 96756
rect 287256 96688 287284 96840
rect 308214 96772 308220 96824
rect 308272 96812 308278 96824
rect 315298 96812 315304 96824
rect 308272 96784 315304 96812
rect 308272 96772 308278 96784
rect 315298 96772 315304 96784
rect 315356 96772 315362 96824
rect 316310 96772 316316 96824
rect 316368 96812 316374 96824
rect 323578 96812 323584 96824
rect 316368 96784 323584 96812
rect 316368 96772 316374 96784
rect 323578 96772 323584 96784
rect 323636 96772 323642 96824
rect 330110 96772 330116 96824
rect 330168 96812 330174 96824
rect 332042 96812 332048 96824
rect 330168 96784 332048 96812
rect 330168 96772 330174 96784
rect 332042 96772 332048 96784
rect 332100 96772 332106 96824
rect 335630 96772 335636 96824
rect 335688 96812 335694 96824
rect 335998 96812 336004 96824
rect 335688 96784 336004 96812
rect 335688 96772 335694 96784
rect 335998 96772 336004 96784
rect 336056 96772 336062 96824
rect 247678 96636 247684 96688
rect 247736 96676 247742 96688
rect 248414 96676 248420 96688
rect 247736 96648 248420 96676
rect 247736 96636 247742 96648
rect 248414 96636 248420 96648
rect 248472 96636 248478 96688
rect 265618 96636 265624 96688
rect 265676 96676 265682 96688
rect 268378 96676 268384 96688
rect 265676 96648 268384 96676
rect 265676 96636 265682 96648
rect 268378 96636 268384 96648
rect 268436 96636 268442 96688
rect 268470 96636 268476 96688
rect 268528 96676 268534 96688
rect 271046 96676 271052 96688
rect 268528 96648 271052 96676
rect 268528 96636 268534 96648
rect 271046 96636 271052 96648
rect 271104 96636 271110 96688
rect 273898 96636 273904 96688
rect 273956 96676 273962 96688
rect 274358 96676 274364 96688
rect 273956 96648 274364 96676
rect 273956 96636 273962 96648
rect 274358 96636 274364 96648
rect 274416 96636 274422 96688
rect 278130 96636 278136 96688
rect 278188 96676 278194 96688
rect 281442 96676 281448 96688
rect 278188 96648 281448 96676
rect 278188 96636 278194 96648
rect 281442 96636 281448 96648
rect 281500 96636 281506 96688
rect 287238 96636 287244 96688
rect 287296 96636 287302 96688
rect 340874 96636 340880 96688
rect 340932 96676 340938 96688
rect 341886 96676 341892 96688
rect 340932 96648 341892 96676
rect 340932 96636 340938 96648
rect 341886 96636 341892 96648
rect 341944 96636 341950 96688
rect 275186 96336 275192 96348
rect 258046 96308 275192 96336
rect 209774 96160 209780 96212
rect 209832 96200 209838 96212
rect 258046 96200 258074 96308
rect 275186 96296 275192 96308
rect 275244 96296 275250 96348
rect 273714 96200 273720 96212
rect 209832 96172 258074 96200
rect 263566 96172 273720 96200
rect 209832 96160 209838 96172
rect 201494 96092 201500 96144
rect 201552 96132 201558 96144
rect 263566 96132 263594 96172
rect 273714 96160 273720 96172
rect 273772 96160 273778 96212
rect 307754 96160 307760 96212
rect 307812 96200 307818 96212
rect 367094 96200 367100 96212
rect 307812 96172 367100 96200
rect 307812 96160 307818 96172
rect 367094 96160 367100 96172
rect 367152 96160 367158 96212
rect 201552 96104 263594 96132
rect 201552 96092 201558 96104
rect 308950 96092 308956 96144
rect 309008 96132 309014 96144
rect 373994 96132 374000 96144
rect 309008 96104 374000 96132
rect 309008 96092 309014 96104
rect 373994 96092 374000 96104
rect 374052 96092 374058 96144
rect 182174 96024 182180 96076
rect 182232 96064 182238 96076
rect 269574 96064 269580 96076
rect 182232 96036 269580 96064
rect 182232 96024 182238 96036
rect 269574 96024 269580 96036
rect 269632 96024 269638 96076
rect 321186 96024 321192 96076
rect 321244 96064 321250 96076
rect 431954 96064 431960 96076
rect 321244 96036 431960 96064
rect 321244 96024 321250 96036
rect 431954 96024 431960 96036
rect 432012 96024 432018 96076
rect 80054 95956 80060 96008
rect 80112 95996 80118 96008
rect 248598 95996 248604 96008
rect 80112 95968 248604 95996
rect 80112 95956 80118 95968
rect 248598 95956 248604 95968
rect 248656 95956 248662 96008
rect 333054 95956 333060 96008
rect 333112 95996 333118 96008
rect 489914 95996 489920 96008
rect 333112 95968 489920 95996
rect 333112 95956 333118 95968
rect 489914 95956 489920 95968
rect 489972 95956 489978 96008
rect 4798 95888 4804 95940
rect 4856 95928 4862 95940
rect 232130 95928 232136 95940
rect 4856 95900 232136 95928
rect 4856 95888 4862 95900
rect 232130 95888 232136 95900
rect 232188 95888 232194 95940
rect 300210 95888 300216 95940
rect 300268 95928 300274 95940
rect 331214 95928 331220 95940
rect 300268 95900 331220 95928
rect 300268 95888 300274 95900
rect 331214 95888 331220 95900
rect 331272 95888 331278 95940
rect 344002 95888 344008 95940
rect 344060 95928 344066 95940
rect 543734 95928 543740 95940
rect 344060 95900 543740 95928
rect 344060 95888 344066 95900
rect 543734 95888 543740 95900
rect 543792 95888 543798 95940
rect 326338 95752 326344 95804
rect 326396 95792 326402 95804
rect 326798 95792 326804 95804
rect 326396 95764 326804 95792
rect 326396 95752 326402 95764
rect 326798 95752 326804 95764
rect 326856 95752 326862 95804
rect 257154 95412 257160 95464
rect 257212 95452 257218 95464
rect 257338 95452 257344 95464
rect 257212 95424 257344 95452
rect 257212 95412 257218 95424
rect 257338 95412 257344 95424
rect 257396 95412 257402 95464
rect 284478 95344 284484 95396
rect 284536 95384 284542 95396
rect 285582 95384 285588 95396
rect 284536 95356 285588 95384
rect 284536 95344 284542 95356
rect 285582 95344 285588 95356
rect 285640 95344 285646 95396
rect 310974 95344 310980 95396
rect 311032 95384 311038 95396
rect 311250 95384 311256 95396
rect 311032 95356 311256 95384
rect 311032 95344 311038 95356
rect 311250 95344 311256 95356
rect 311308 95344 311314 95396
rect 268194 94800 268200 94852
rect 268252 94840 268258 94852
rect 268654 94840 268660 94852
rect 268252 94812 268660 94840
rect 268252 94800 268258 94812
rect 268654 94800 268660 94812
rect 268712 94800 268718 94852
rect 264146 94732 264152 94784
rect 264204 94772 264210 94784
rect 264514 94772 264520 94784
rect 264204 94744 264520 94772
rect 264204 94732 264210 94744
rect 264514 94732 264520 94744
rect 264572 94732 264578 94784
rect 267918 94732 267924 94784
rect 267976 94772 267982 94784
rect 268562 94772 268568 94784
rect 267976 94744 268568 94772
rect 267976 94732 267982 94744
rect 268562 94732 268568 94744
rect 268620 94732 268626 94784
rect 305362 94732 305368 94784
rect 305420 94772 305426 94784
rect 356054 94772 356060 94784
rect 305420 94744 356060 94772
rect 305420 94732 305426 94744
rect 356054 94732 356060 94744
rect 356112 94732 356118 94784
rect 227714 94664 227720 94716
rect 227772 94704 227778 94716
rect 279050 94704 279056 94716
rect 227772 94676 279056 94704
rect 227772 94664 227778 94676
rect 279050 94664 279056 94676
rect 279108 94664 279114 94716
rect 306926 94664 306932 94716
rect 306984 94704 306990 94716
rect 364334 94704 364340 94716
rect 306984 94676 364340 94704
rect 306984 94664 306990 94676
rect 364334 94664 364340 94676
rect 364392 94664 364398 94716
rect 195974 94596 195980 94648
rect 196032 94636 196038 94648
rect 270494 94636 270500 94648
rect 196032 94608 270500 94636
rect 196032 94596 196038 94608
rect 270494 94596 270500 94608
rect 270552 94596 270558 94648
rect 311618 94596 311624 94648
rect 311676 94636 311682 94648
rect 386414 94636 386420 94648
rect 311676 94608 386420 94636
rect 311676 94596 311682 94608
rect 386414 94596 386420 94608
rect 386472 94596 386478 94648
rect 125594 94528 125600 94580
rect 125652 94568 125658 94580
rect 257890 94568 257896 94580
rect 125652 94540 257896 94568
rect 125652 94528 125658 94540
rect 257890 94528 257896 94540
rect 257948 94528 257954 94580
rect 263962 94528 263968 94580
rect 264020 94568 264026 94580
rect 264514 94568 264520 94580
rect 264020 94540 264520 94568
rect 264020 94528 264026 94540
rect 264514 94528 264520 94540
rect 264572 94528 264578 94580
rect 266722 94528 266728 94580
rect 266780 94568 266786 94580
rect 267090 94568 267096 94580
rect 266780 94540 267096 94568
rect 266780 94528 266786 94540
rect 267090 94528 267096 94540
rect 267148 94528 267154 94580
rect 269114 94528 269120 94580
rect 269172 94568 269178 94580
rect 270126 94568 270132 94580
rect 269172 94540 270132 94568
rect 269172 94528 269178 94540
rect 270126 94528 270132 94540
rect 270184 94528 270190 94580
rect 270862 94528 270868 94580
rect 270920 94568 270926 94580
rect 271598 94568 271604 94580
rect 270920 94540 271604 94568
rect 270920 94528 270926 94540
rect 271598 94528 271604 94540
rect 271656 94528 271662 94580
rect 272058 94528 272064 94580
rect 272116 94568 272122 94580
rect 272702 94568 272708 94580
rect 272116 94540 272708 94568
rect 272116 94528 272122 94540
rect 272702 94528 272708 94540
rect 272760 94528 272766 94580
rect 333790 94528 333796 94580
rect 333848 94568 333854 94580
rect 494054 94568 494060 94580
rect 333848 94540 494060 94568
rect 333848 94528 333854 94540
rect 494054 94528 494060 94540
rect 494112 94528 494118 94580
rect 60734 94460 60740 94512
rect 60792 94500 60798 94512
rect 242986 94500 242992 94512
rect 60792 94472 242992 94500
rect 60792 94460 60798 94472
rect 242986 94460 242992 94472
rect 243044 94460 243050 94512
rect 246298 94460 246304 94512
rect 246356 94500 246362 94512
rect 246666 94500 246672 94512
rect 246356 94472 246672 94500
rect 246356 94460 246362 94472
rect 246666 94460 246672 94472
rect 246724 94460 246730 94512
rect 247494 94460 247500 94512
rect 247552 94500 247558 94512
rect 247954 94500 247960 94512
rect 247552 94472 247960 94500
rect 247552 94460 247558 94472
rect 247954 94460 247960 94472
rect 248012 94460 248018 94512
rect 248690 94460 248696 94512
rect 248748 94500 248754 94512
rect 248966 94500 248972 94512
rect 248748 94472 248972 94500
rect 248748 94460 248754 94472
rect 248966 94460 248972 94472
rect 249024 94460 249030 94512
rect 250162 94460 250168 94512
rect 250220 94500 250226 94512
rect 250438 94500 250444 94512
rect 250220 94472 250444 94500
rect 250220 94460 250226 94472
rect 250438 94460 250444 94472
rect 250496 94460 250502 94512
rect 251358 94460 251364 94512
rect 251416 94500 251422 94512
rect 252094 94500 252100 94512
rect 251416 94472 252100 94500
rect 251416 94460 251422 94472
rect 252094 94460 252100 94472
rect 252152 94460 252158 94512
rect 252554 94460 252560 94512
rect 252612 94500 252618 94512
rect 252830 94500 252836 94512
rect 252612 94472 252836 94500
rect 252612 94460 252618 94472
rect 252830 94460 252836 94472
rect 252888 94460 252894 94512
rect 267826 94460 267832 94512
rect 267884 94500 267890 94512
rect 268654 94500 268660 94512
rect 267884 94472 268660 94500
rect 267884 94460 267890 94472
rect 268654 94460 268660 94472
rect 268712 94460 268718 94512
rect 270586 94460 270592 94512
rect 270644 94500 270650 94512
rect 271322 94500 271328 94512
rect 270644 94472 271328 94500
rect 270644 94460 270650 94472
rect 271322 94460 271328 94472
rect 271380 94460 271386 94512
rect 346946 94460 346952 94512
rect 347004 94500 347010 94512
rect 557534 94500 557540 94512
rect 347004 94472 557540 94500
rect 347004 94460 347010 94472
rect 557534 94460 557540 94472
rect 557592 94460 557598 94512
rect 247218 94392 247224 94444
rect 247276 94432 247282 94444
rect 247862 94432 247868 94444
rect 247276 94404 247868 94432
rect 247276 94392 247282 94404
rect 247862 94392 247868 94404
rect 247920 94392 247926 94444
rect 248966 94324 248972 94376
rect 249024 94364 249030 94376
rect 249426 94364 249432 94376
rect 249024 94336 249432 94364
rect 249024 94324 249030 94336
rect 249426 94324 249432 94336
rect 249484 94324 249490 94376
rect 250438 94324 250444 94376
rect 250496 94364 250502 94376
rect 250898 94364 250904 94376
rect 250496 94336 250904 94364
rect 250496 94324 250502 94336
rect 250898 94324 250904 94336
rect 250956 94324 250962 94376
rect 270586 94324 270592 94376
rect 270644 94364 270650 94376
rect 271506 94364 271512 94376
rect 270644 94336 271512 94364
rect 270644 94324 270650 94336
rect 271506 94324 271512 94336
rect 271564 94324 271570 94376
rect 304626 93372 304632 93424
rect 304684 93412 304690 93424
rect 351914 93412 351920 93424
rect 304684 93384 351920 93412
rect 304684 93372 304690 93384
rect 351914 93372 351920 93384
rect 351972 93372 351978 93424
rect 200114 93304 200120 93356
rect 200172 93344 200178 93356
rect 273254 93344 273260 93356
rect 200172 93316 273260 93344
rect 200172 93304 200178 93316
rect 273254 93304 273260 93316
rect 273312 93304 273318 93356
rect 332134 93304 332140 93356
rect 332192 93344 332198 93356
rect 387794 93344 387800 93356
rect 332192 93316 387800 93344
rect 332192 93304 332198 93316
rect 387794 93304 387800 93316
rect 387852 93304 387858 93356
rect 193214 93236 193220 93288
rect 193272 93276 193278 93288
rect 271966 93276 271972 93288
rect 193272 93248 271972 93276
rect 193272 93236 193278 93248
rect 271966 93236 271972 93248
rect 272024 93236 272030 93288
rect 326522 93236 326528 93288
rect 326580 93276 326586 93288
rect 458174 93276 458180 93288
rect 326580 93248 458180 93276
rect 326580 93236 326586 93248
rect 458174 93236 458180 93248
rect 458232 93236 458238 93288
rect 160094 93168 160100 93220
rect 160152 93208 160158 93220
rect 257430 93208 257436 93220
rect 160152 93180 257436 93208
rect 160152 93168 160158 93180
rect 257430 93168 257436 93180
rect 257488 93168 257494 93220
rect 336182 93168 336188 93220
rect 336240 93208 336246 93220
rect 498194 93208 498200 93220
rect 336240 93180 498200 93208
rect 336240 93168 336246 93180
rect 498194 93168 498200 93180
rect 498252 93168 498258 93220
rect 71774 93100 71780 93152
rect 71832 93140 71838 93152
rect 246758 93140 246764 93152
rect 71832 93112 246764 93140
rect 71832 93100 71838 93112
rect 246758 93100 246764 93112
rect 246816 93100 246822 93152
rect 351086 93100 351092 93152
rect 351144 93140 351150 93152
rect 578234 93140 578240 93152
rect 351144 93112 578240 93140
rect 351144 93100 351150 93112
rect 578234 93100 578240 93112
rect 578292 93100 578298 93152
rect 215294 92012 215300 92064
rect 215352 92052 215358 92064
rect 276382 92052 276388 92064
rect 215352 92024 276388 92052
rect 215352 92012 215358 92024
rect 276382 92012 276388 92024
rect 276440 92012 276446 92064
rect 207014 91944 207020 91996
rect 207072 91984 207078 91996
rect 274634 91984 274640 91996
rect 207072 91956 274640 91984
rect 207072 91944 207078 91956
rect 274634 91944 274640 91956
rect 274692 91944 274698 91996
rect 305914 91944 305920 91996
rect 305972 91984 305978 91996
rect 358814 91984 358820 91996
rect 305972 91956 358820 91984
rect 305972 91944 305978 91956
rect 358814 91944 358820 91956
rect 358872 91944 358878 91996
rect 164234 91876 164240 91928
rect 164292 91916 164298 91928
rect 265894 91916 265900 91928
rect 164292 91888 265900 91916
rect 164292 91876 164298 91888
rect 265894 91876 265900 91888
rect 265952 91876 265958 91928
rect 312630 91876 312636 91928
rect 312688 91916 312694 91928
rect 390554 91916 390560 91928
rect 312688 91888 390560 91916
rect 312688 91876 312694 91888
rect 390554 91876 390560 91888
rect 390612 91876 390618 91928
rect 113174 91808 113180 91860
rect 113232 91848 113238 91860
rect 255406 91848 255412 91860
rect 113232 91820 255412 91848
rect 113232 91808 113238 91820
rect 255406 91808 255412 91820
rect 255464 91808 255470 91860
rect 336734 91808 336740 91860
rect 336792 91848 336798 91860
rect 507854 91848 507860 91860
rect 336792 91820 507860 91848
rect 336792 91808 336798 91820
rect 507854 91808 507860 91820
rect 507912 91808 507918 91860
rect 46934 91740 46940 91792
rect 46992 91780 46998 91792
rect 241882 91780 241888 91792
rect 46992 91752 241888 91780
rect 46992 91740 46998 91752
rect 241882 91740 241888 91752
rect 241940 91740 241946 91792
rect 344278 91740 344284 91792
rect 344336 91780 344342 91792
rect 545114 91780 545120 91792
rect 344336 91752 545120 91780
rect 344336 91740 344342 91752
rect 545114 91740 545120 91752
rect 545172 91740 545178 91792
rect 213914 90516 213920 90568
rect 213972 90556 213978 90568
rect 275462 90556 275468 90568
rect 213972 90528 275468 90556
rect 213972 90516 213978 90528
rect 275462 90516 275468 90528
rect 275520 90516 275526 90568
rect 306834 90516 306840 90568
rect 306892 90556 306898 90568
rect 362954 90556 362960 90568
rect 306892 90528 362960 90556
rect 306892 90516 306898 90528
rect 362954 90516 362960 90528
rect 363012 90516 363018 90568
rect 171134 90448 171140 90500
rect 171192 90488 171198 90500
rect 265434 90488 265440 90500
rect 171192 90460 265440 90488
rect 171192 90448 171198 90460
rect 265434 90448 265440 90460
rect 265492 90448 265498 90500
rect 313366 90448 313372 90500
rect 313424 90488 313430 90500
rect 394694 90488 394700 90500
rect 313424 90460 394700 90488
rect 313424 90448 313430 90460
rect 394694 90448 394700 90460
rect 394752 90448 394758 90500
rect 151814 90380 151820 90432
rect 151872 90420 151878 90432
rect 263042 90420 263048 90432
rect 151872 90392 263048 90420
rect 151872 90380 151878 90392
rect 263042 90380 263048 90392
rect 263100 90380 263106 90432
rect 337470 90380 337476 90432
rect 337528 90420 337534 90432
rect 511994 90420 512000 90432
rect 337528 90392 512000 90420
rect 337528 90380 337534 90392
rect 511994 90380 512000 90392
rect 512052 90380 512058 90432
rect 26234 90312 26240 90364
rect 26292 90352 26298 90364
rect 237466 90352 237472 90364
rect 26292 90324 237472 90352
rect 26292 90312 26298 90324
rect 237466 90312 237472 90324
rect 237524 90312 237530 90364
rect 347958 90312 347964 90364
rect 348016 90352 348022 90364
rect 563054 90352 563060 90364
rect 348016 90324 563060 90352
rect 348016 90312 348022 90324
rect 563054 90312 563060 90324
rect 563112 90312 563118 90364
rect 265158 90108 265164 90160
rect 265216 90148 265222 90160
rect 265526 90148 265532 90160
rect 265216 90120 265532 90148
rect 265216 90108 265222 90120
rect 265526 90108 265532 90120
rect 265584 90108 265590 90160
rect 220814 89156 220820 89208
rect 220872 89196 220878 89208
rect 277670 89196 277676 89208
rect 220872 89168 277676 89196
rect 220872 89156 220878 89168
rect 277670 89156 277676 89168
rect 277728 89156 277734 89208
rect 315298 89156 315304 89208
rect 315356 89196 315362 89208
rect 369854 89196 369860 89208
rect 315356 89168 369860 89196
rect 315356 89156 315362 89168
rect 369854 89156 369860 89168
rect 369912 89156 369918 89208
rect 175274 89088 175280 89140
rect 175332 89128 175338 89140
rect 268102 89128 268108 89140
rect 175332 89100 268108 89128
rect 175332 89088 175338 89100
rect 268102 89088 268108 89100
rect 268160 89088 268166 89140
rect 319162 89088 319168 89140
rect 319220 89128 319226 89140
rect 423674 89128 423680 89140
rect 319220 89100 423680 89128
rect 319220 89088 319226 89100
rect 423674 89088 423680 89100
rect 423732 89088 423738 89140
rect 147674 89020 147680 89072
rect 147732 89060 147738 89072
rect 262490 89060 262496 89072
rect 147732 89032 262496 89060
rect 147732 89020 147738 89032
rect 262490 89020 262496 89032
rect 262548 89020 262554 89072
rect 325142 89020 325148 89072
rect 325200 89060 325206 89072
rect 452654 89060 452660 89072
rect 325200 89032 452660 89060
rect 325200 89020 325206 89032
rect 452654 89020 452660 89032
rect 452712 89020 452718 89072
rect 16574 88952 16580 89004
rect 16632 88992 16638 89004
rect 234614 88992 234620 89004
rect 16632 88964 234620 88992
rect 16632 88952 16638 88964
rect 234614 88952 234620 88964
rect 234672 88952 234678 89004
rect 338942 88952 338948 89004
rect 339000 88992 339006 89004
rect 518894 88992 518900 89004
rect 339000 88964 518900 88992
rect 339000 88952 339006 88964
rect 518894 88952 518900 88964
rect 518952 88952 518958 89004
rect 230474 87796 230480 87848
rect 230532 87836 230538 87848
rect 279878 87836 279884 87848
rect 230532 87808 279884 87836
rect 230532 87796 230538 87808
rect 279878 87796 279884 87808
rect 279936 87796 279942 87848
rect 309686 87796 309692 87848
rect 309744 87836 309750 87848
rect 376754 87836 376760 87848
rect 309744 87808 376760 87836
rect 309744 87796 309750 87808
rect 376754 87796 376760 87808
rect 376812 87796 376818 87848
rect 178034 87728 178040 87780
rect 178092 87768 178098 87780
rect 268194 87768 268200 87780
rect 178092 87740 268200 87768
rect 178092 87728 178098 87740
rect 268194 87728 268200 87740
rect 268252 87728 268258 87780
rect 322658 87728 322664 87780
rect 322716 87768 322722 87780
rect 440326 87768 440332 87780
rect 322716 87740 440332 87768
rect 322716 87728 322722 87740
rect 440326 87728 440332 87740
rect 440384 87728 440390 87780
rect 139394 87660 139400 87712
rect 139452 87700 139458 87712
rect 260834 87700 260840 87712
rect 139452 87672 260840 87700
rect 139452 87660 139458 87672
rect 260834 87660 260840 87672
rect 260892 87660 260898 87712
rect 330386 87660 330392 87712
rect 330444 87700 330450 87712
rect 477494 87700 477500 87712
rect 330444 87672 477500 87700
rect 330444 87660 330450 87672
rect 477494 87660 477500 87672
rect 477552 87660 477558 87712
rect 103514 87592 103520 87644
rect 103572 87632 103578 87644
rect 253474 87632 253480 87644
rect 103572 87604 253480 87632
rect 103572 87592 103578 87604
rect 253474 87592 253480 87604
rect 253532 87592 253538 87644
rect 267734 87592 267740 87644
rect 267792 87632 267798 87644
rect 287238 87632 287244 87644
rect 267792 87604 287244 87632
rect 267792 87592 267798 87604
rect 287238 87592 287244 87604
rect 287296 87592 287302 87644
rect 339678 87592 339684 87644
rect 339736 87632 339742 87644
rect 523034 87632 523040 87644
rect 339736 87604 523040 87632
rect 339736 87592 339742 87604
rect 523034 87592 523040 87604
rect 523092 87592 523098 87644
rect 354490 86912 354496 86964
rect 354548 86952 354554 86964
rect 580166 86952 580172 86964
rect 354548 86924 580172 86952
rect 354548 86912 354554 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 219434 86436 219440 86488
rect 219492 86476 219498 86488
rect 276198 86476 276204 86488
rect 219492 86448 276204 86476
rect 219492 86436 219498 86448
rect 276198 86436 276204 86448
rect 276256 86436 276262 86488
rect 184934 86368 184940 86420
rect 184992 86408 184998 86420
rect 270310 86408 270316 86420
rect 184992 86380 270316 86408
rect 184992 86368 184998 86380
rect 270310 86368 270316 86380
rect 270368 86368 270374 86420
rect 306650 86368 306656 86420
rect 306708 86408 306714 86420
rect 365714 86408 365720 86420
rect 306708 86380 365720 86408
rect 306708 86368 306714 86380
rect 365714 86368 365720 86380
rect 365772 86368 365778 86420
rect 146294 86300 146300 86352
rect 146352 86340 146358 86352
rect 260190 86340 260196 86352
rect 146352 86312 260196 86340
rect 146352 86300 146358 86312
rect 260190 86300 260196 86312
rect 260248 86300 260254 86352
rect 323578 86300 323584 86352
rect 323636 86340 323642 86352
rect 408494 86340 408500 86352
rect 323636 86312 408500 86340
rect 323636 86300 323642 86312
rect 408494 86300 408500 86312
rect 408552 86300 408558 86352
rect 20714 86232 20720 86284
rect 20772 86272 20778 86284
rect 233878 86272 233884 86284
rect 20772 86244 233884 86272
rect 20772 86232 20778 86244
rect 233878 86232 233884 86244
rect 233936 86232 233942 86284
rect 316494 86232 316500 86284
rect 316552 86272 316558 86284
rect 409874 86272 409880 86284
rect 316552 86244 409880 86272
rect 316552 86232 316558 86244
rect 409874 86232 409880 86244
rect 409932 86232 409938 86284
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 230106 85524 230112 85536
rect 3384 85496 230112 85524
rect 3384 85484 3390 85496
rect 230106 85484 230112 85496
rect 230164 85484 230170 85536
rect 308030 85008 308036 85060
rect 308088 85048 308094 85060
rect 368474 85048 368480 85060
rect 308088 85020 368480 85048
rect 308088 85008 308094 85020
rect 368474 85008 368480 85020
rect 368532 85008 368538 85060
rect 218054 84940 218060 84992
rect 218112 84980 218118 84992
rect 276934 84980 276940 84992
rect 218112 84952 276940 84980
rect 218112 84940 218118 84952
rect 276934 84940 276940 84952
rect 276992 84940 276998 84992
rect 311066 84940 311072 84992
rect 311124 84980 311130 84992
rect 383654 84980 383660 84992
rect 311124 84952 383660 84980
rect 311124 84940 311130 84952
rect 383654 84940 383660 84952
rect 383712 84940 383718 84992
rect 202874 84872 202880 84924
rect 202932 84912 202938 84924
rect 273806 84912 273812 84924
rect 202932 84884 273812 84912
rect 202932 84872 202938 84884
rect 273806 84872 273812 84884
rect 273864 84872 273870 84924
rect 340230 84872 340236 84924
rect 340288 84912 340294 84924
rect 525794 84912 525800 84924
rect 340288 84884 525800 84912
rect 340288 84872 340294 84884
rect 525794 84872 525800 84884
rect 525852 84872 525858 84924
rect 107654 84804 107660 84856
rect 107712 84844 107718 84856
rect 254302 84844 254308 84856
rect 107712 84816 254308 84844
rect 107712 84804 107718 84816
rect 254302 84804 254308 84816
rect 254360 84804 254366 84856
rect 294598 84804 294604 84856
rect 294656 84844 294662 84856
rect 303614 84844 303620 84856
rect 294656 84816 303620 84844
rect 294656 84804 294662 84816
rect 303614 84804 303620 84816
rect 303672 84804 303678 84856
rect 347774 84804 347780 84856
rect 347832 84844 347838 84856
rect 565814 84844 565820 84856
rect 347832 84816 565820 84844
rect 347832 84804 347838 84816
rect 565814 84804 565820 84816
rect 565872 84804 565878 84856
rect 310054 83648 310060 83700
rect 310112 83688 310118 83700
rect 380894 83688 380900 83700
rect 310112 83660 380900 83688
rect 310112 83648 310118 83660
rect 380894 83648 380900 83660
rect 380952 83648 380958 83700
rect 189074 83580 189080 83632
rect 189132 83620 189138 83632
rect 268470 83620 268476 83632
rect 189132 83592 268476 83620
rect 189132 83580 189138 83592
rect 268470 83580 268476 83592
rect 268528 83580 268534 83632
rect 355502 83580 355508 83632
rect 355560 83620 355566 83632
rect 480254 83620 480260 83632
rect 355560 83592 480260 83620
rect 355560 83580 355566 83592
rect 480254 83580 480260 83592
rect 480312 83580 480318 83632
rect 126974 83512 126980 83564
rect 127032 83552 127038 83564
rect 258166 83552 258172 83564
rect 127032 83524 258172 83552
rect 127032 83512 127038 83524
rect 258166 83512 258172 83524
rect 258224 83512 258230 83564
rect 327718 83512 327724 83564
rect 327776 83552 327782 83564
rect 455414 83552 455420 83564
rect 327776 83524 455420 83552
rect 327776 83512 327782 83524
rect 455414 83512 455420 83524
rect 455472 83512 455478 83564
rect 85574 83444 85580 83496
rect 85632 83484 85638 83496
rect 249794 83484 249800 83496
rect 85632 83456 249800 83484
rect 85632 83444 85638 83456
rect 249794 83444 249800 83456
rect 249852 83444 249858 83496
rect 267826 83444 267832 83496
rect 267884 83484 267890 83496
rect 287422 83484 287428 83496
rect 267884 83456 287428 83484
rect 267884 83444 267890 83456
rect 287422 83444 287428 83456
rect 287480 83444 287486 83496
rect 349522 83444 349528 83496
rect 349580 83484 349586 83496
rect 571334 83484 571340 83496
rect 349580 83456 571340 83484
rect 349580 83444 349586 83456
rect 571334 83444 571340 83456
rect 571392 83444 571398 83496
rect 193306 82220 193312 82272
rect 193364 82260 193370 82272
rect 270862 82260 270868 82272
rect 193364 82232 270868 82260
rect 193364 82220 193370 82232
rect 270862 82220 270868 82232
rect 270920 82220 270926 82272
rect 312078 82220 312084 82272
rect 312136 82260 312142 82272
rect 389174 82260 389180 82272
rect 312136 82232 389180 82260
rect 312136 82220 312142 82232
rect 389174 82220 389180 82232
rect 389232 82220 389238 82272
rect 129734 82152 129740 82204
rect 129792 82192 129798 82204
rect 258718 82192 258724 82204
rect 129792 82164 258724 82192
rect 129792 82152 129798 82164
rect 258718 82152 258724 82164
rect 258776 82152 258782 82204
rect 333330 82152 333336 82204
rect 333388 82192 333394 82204
rect 412634 82192 412640 82204
rect 333388 82164 412640 82192
rect 333388 82152 333394 82164
rect 412634 82152 412640 82164
rect 412692 82152 412698 82204
rect 89714 82084 89720 82136
rect 89772 82124 89778 82136
rect 250162 82124 250168 82136
rect 89772 82096 250168 82124
rect 89772 82084 89778 82096
rect 250162 82084 250168 82096
rect 250220 82084 250226 82136
rect 302326 82084 302332 82136
rect 302384 82124 302390 82136
rect 340874 82124 340880 82136
rect 302384 82096 340880 82124
rect 302384 82084 302390 82096
rect 340874 82084 340880 82096
rect 340932 82084 340938 82136
rect 340966 82084 340972 82136
rect 341024 82124 341030 82136
rect 529934 82124 529940 82136
rect 341024 82096 529940 82124
rect 341024 82084 341030 82096
rect 529934 82084 529940 82096
rect 529992 82084 529998 82136
rect 308306 80860 308312 80912
rect 308364 80900 308370 80912
rect 371234 80900 371240 80912
rect 308364 80872 371240 80900
rect 308364 80860 308370 80872
rect 371234 80860 371240 80872
rect 371292 80860 371298 80912
rect 211154 80792 211160 80844
rect 211212 80832 211218 80844
rect 275554 80832 275560 80844
rect 211212 80804 275560 80832
rect 211212 80792 211218 80804
rect 275554 80792 275560 80804
rect 275612 80792 275618 80844
rect 314010 80792 314016 80844
rect 314068 80832 314074 80844
rect 398834 80832 398840 80844
rect 314068 80804 398840 80832
rect 314068 80792 314074 80804
rect 398834 80792 398840 80804
rect 398892 80792 398898 80844
rect 128354 80724 128360 80776
rect 128412 80764 128418 80776
rect 257338 80764 257344 80776
rect 128412 80736 257344 80764
rect 128412 80724 128418 80736
rect 257338 80724 257344 80736
rect 257396 80724 257402 80776
rect 326614 80724 326620 80776
rect 326672 80764 326678 80776
rect 459554 80764 459560 80776
rect 326672 80736 459560 80764
rect 326672 80724 326678 80736
rect 459554 80724 459560 80736
rect 459612 80724 459618 80776
rect 78674 80656 78680 80708
rect 78732 80696 78738 80708
rect 247678 80696 247684 80708
rect 78732 80668 247684 80696
rect 78732 80656 78738 80668
rect 247678 80656 247684 80668
rect 247736 80656 247742 80708
rect 256786 80656 256792 80708
rect 256844 80696 256850 80708
rect 284754 80696 284760 80708
rect 256844 80668 284760 80696
rect 256844 80656 256850 80668
rect 284754 80656 284760 80668
rect 284812 80656 284818 80708
rect 342438 80656 342444 80708
rect 342496 80696 342502 80708
rect 536834 80696 536840 80708
rect 342496 80668 536840 80696
rect 342496 80656 342502 80668
rect 536834 80656 536840 80668
rect 536892 80656 536898 80708
rect 224954 79500 224960 79552
rect 225012 79540 225018 79552
rect 278222 79540 278228 79552
rect 225012 79512 278228 79540
rect 225012 79500 225018 79512
rect 278222 79500 278228 79512
rect 278280 79500 278286 79552
rect 150434 79432 150440 79484
rect 150492 79472 150498 79484
rect 261478 79472 261484 79484
rect 150492 79444 261484 79472
rect 150492 79432 150498 79444
rect 261478 79432 261484 79444
rect 261536 79432 261542 79484
rect 312446 79432 312452 79484
rect 312504 79472 312510 79484
rect 391934 79472 391940 79484
rect 312504 79444 391940 79472
rect 312504 79432 312510 79444
rect 391934 79432 391940 79444
rect 391992 79432 391998 79484
rect 53834 79364 53840 79416
rect 53892 79404 53898 79416
rect 243262 79404 243268 79416
rect 53892 79376 243268 79404
rect 53892 79364 53898 79376
rect 243262 79364 243268 79376
rect 243320 79364 243326 79416
rect 317690 79364 317696 79416
rect 317748 79404 317754 79416
rect 415394 79404 415400 79416
rect 317748 79376 415400 79404
rect 317748 79364 317754 79376
rect 415394 79364 415400 79376
rect 415452 79364 415458 79416
rect 13814 79296 13820 79348
rect 13872 79336 13878 79348
rect 234890 79336 234896 79348
rect 13872 79308 234896 79336
rect 13872 79296 13878 79308
rect 234890 79296 234896 79308
rect 234948 79296 234954 79348
rect 343174 79296 343180 79348
rect 343232 79336 343238 79348
rect 539594 79336 539600 79348
rect 343232 79308 539600 79336
rect 343232 79296 343238 79308
rect 539594 79296 539600 79308
rect 539652 79296 539658 79348
rect 197354 78072 197360 78124
rect 197412 78112 197418 78124
rect 272058 78112 272064 78124
rect 197412 78084 272064 78112
rect 197412 78072 197418 78084
rect 272058 78072 272064 78084
rect 272116 78072 272122 78124
rect 316586 78072 316592 78124
rect 316644 78112 316650 78124
rect 414014 78112 414020 78124
rect 316644 78084 414020 78112
rect 316644 78072 316650 78084
rect 414014 78072 414020 78084
rect 414072 78072 414078 78124
rect 132494 78004 132500 78056
rect 132552 78044 132558 78056
rect 255958 78044 255964 78056
rect 132552 78016 255964 78044
rect 132552 78004 132558 78016
rect 255958 78004 255964 78016
rect 256016 78004 256022 78056
rect 320542 78004 320548 78056
rect 320600 78044 320606 78056
rect 430574 78044 430580 78056
rect 320600 78016 430580 78044
rect 320600 78004 320606 78016
rect 430574 78004 430580 78016
rect 430632 78004 430638 78056
rect 100754 77936 100760 77988
rect 100812 77976 100818 77988
rect 252646 77976 252652 77988
rect 100812 77948 252652 77976
rect 100812 77936 100818 77948
rect 252646 77936 252652 77948
rect 252704 77936 252710 77988
rect 344094 77936 344100 77988
rect 344152 77976 344158 77988
rect 547874 77976 547880 77988
rect 344152 77948 547880 77976
rect 344152 77936 344158 77948
rect 547874 77936 547880 77948
rect 547932 77936 547938 77988
rect 231854 76712 231860 76764
rect 231912 76752 231918 76764
rect 279694 76752 279700 76764
rect 231912 76724 279700 76752
rect 231912 76712 231918 76724
rect 279694 76712 279700 76724
rect 279752 76712 279758 76764
rect 168374 76644 168380 76696
rect 168432 76684 168438 76696
rect 266814 76684 266820 76696
rect 168432 76656 266820 76684
rect 168432 76644 168438 76656
rect 266814 76644 266820 76656
rect 266872 76644 266878 76696
rect 324314 76644 324320 76696
rect 324372 76684 324378 76696
rect 448514 76684 448520 76696
rect 324372 76656 448520 76684
rect 324372 76644 324378 76656
rect 448514 76644 448520 76656
rect 448572 76644 448578 76696
rect 41414 76576 41420 76628
rect 41472 76616 41478 76628
rect 240410 76616 240416 76628
rect 41472 76588 240416 76616
rect 41472 76576 41478 76588
rect 240410 76576 240416 76588
rect 240468 76576 240474 76628
rect 331950 76576 331956 76628
rect 332008 76616 332014 76628
rect 485774 76616 485780 76628
rect 332008 76588 485780 76616
rect 332008 76576 332014 76588
rect 485774 76576 485780 76588
rect 485832 76576 485838 76628
rect 7558 76508 7564 76560
rect 7616 76548 7622 76560
rect 232222 76548 232228 76560
rect 7616 76520 232228 76548
rect 7616 76508 7622 76520
rect 232222 76508 232228 76520
rect 232280 76508 232286 76560
rect 346026 76508 346032 76560
rect 346084 76548 346090 76560
rect 554774 76548 554780 76560
rect 346084 76520 554780 76548
rect 346084 76508 346090 76520
rect 554774 76508 554780 76520
rect 554832 76508 554838 76560
rect 304442 75352 304448 75404
rect 304500 75392 304506 75404
rect 347774 75392 347780 75404
rect 304500 75364 347780 75392
rect 304500 75352 304506 75364
rect 347774 75352 347780 75364
rect 347832 75352 347838 75404
rect 173894 75284 173900 75336
rect 173952 75324 173958 75336
rect 268654 75324 268660 75336
rect 173952 75296 268660 75324
rect 173952 75284 173958 75296
rect 268654 75284 268660 75296
rect 268712 75284 268718 75336
rect 312262 75284 312268 75336
rect 312320 75324 312326 75336
rect 390646 75324 390652 75336
rect 312320 75296 390652 75324
rect 312320 75284 312326 75296
rect 390646 75284 390652 75296
rect 390704 75284 390710 75336
rect 135254 75216 135260 75268
rect 135312 75256 135318 75268
rect 260006 75256 260012 75268
rect 135312 75228 260012 75256
rect 135312 75216 135318 75228
rect 260006 75216 260012 75228
rect 260064 75216 260070 75268
rect 330478 75216 330484 75268
rect 330536 75256 330542 75268
rect 481634 75256 481640 75268
rect 330536 75228 481640 75256
rect 330536 75216 330542 75228
rect 481634 75216 481640 75228
rect 481692 75216 481698 75268
rect 40034 75148 40040 75200
rect 40092 75188 40098 75200
rect 239398 75188 239404 75200
rect 40092 75160 239404 75188
rect 40092 75148 40098 75160
rect 239398 75148 239404 75160
rect 239456 75148 239462 75200
rect 347498 75148 347504 75200
rect 347556 75188 347562 75200
rect 561674 75188 561680 75200
rect 347556 75160 561680 75188
rect 347556 75148 347562 75160
rect 561674 75148 561680 75160
rect 561732 75148 561738 75200
rect 305454 73992 305460 74044
rect 305512 74032 305518 74044
rect 357434 74032 357440 74044
rect 305512 74004 357440 74032
rect 305512 73992 305518 74004
rect 357434 73992 357440 74004
rect 357492 73992 357498 74044
rect 180794 73924 180800 73976
rect 180852 73964 180858 73976
rect 269390 73964 269396 73976
rect 180852 73936 269396 73964
rect 180852 73924 180858 73936
rect 269390 73924 269396 73936
rect 269448 73924 269454 73976
rect 309778 73924 309784 73976
rect 309836 73964 309842 73976
rect 378134 73964 378140 73976
rect 309836 73936 378140 73964
rect 309836 73924 309842 73936
rect 378134 73924 378140 73936
rect 378192 73924 378198 73976
rect 143534 73856 143540 73908
rect 143592 73896 143598 73908
rect 261110 73896 261116 73908
rect 143592 73868 261116 73896
rect 143592 73856 143598 73868
rect 261110 73856 261116 73868
rect 261168 73856 261174 73908
rect 323026 73856 323032 73908
rect 323084 73896 323090 73908
rect 441614 73896 441620 73908
rect 323084 73868 441620 73896
rect 323084 73856 323090 73868
rect 441614 73856 441620 73868
rect 441672 73856 441678 73908
rect 35894 73788 35900 73840
rect 35952 73828 35958 73840
rect 239490 73828 239496 73840
rect 35952 73800 239496 73828
rect 35952 73788 35958 73800
rect 239490 73788 239496 73800
rect 239548 73788 239554 73840
rect 352742 73788 352748 73840
rect 352800 73828 352806 73840
rect 564526 73828 564532 73840
rect 352800 73800 564532 73828
rect 352800 73788 352806 73800
rect 564526 73788 564532 73800
rect 564584 73788 564590 73840
rect 354398 73108 354404 73160
rect 354456 73148 354462 73160
rect 580166 73148 580172 73160
rect 354456 73120 580172 73148
rect 354456 73108 354462 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 198734 72564 198740 72616
rect 198792 72604 198798 72616
rect 272794 72604 272800 72616
rect 198792 72576 272800 72604
rect 198792 72564 198798 72576
rect 272794 72564 272800 72576
rect 272852 72564 272858 72616
rect 305638 72564 305644 72616
rect 305696 72604 305702 72616
rect 360194 72604 360200 72616
rect 305696 72576 360200 72604
rect 305696 72564 305702 72576
rect 360194 72564 360200 72576
rect 360252 72564 360258 72616
rect 153194 72496 153200 72548
rect 153252 72536 153258 72548
rect 263594 72536 263600 72548
rect 153252 72508 263600 72536
rect 153252 72496 153258 72508
rect 263594 72496 263600 72508
rect 263652 72496 263658 72548
rect 310974 72496 310980 72548
rect 311032 72536 311038 72548
rect 385034 72536 385040 72548
rect 311032 72508 385040 72536
rect 311032 72496 311038 72508
rect 385034 72496 385040 72508
rect 385092 72496 385098 72548
rect 28994 72428 29000 72480
rect 29052 72468 29058 72480
rect 237742 72468 237748 72480
rect 29052 72440 237748 72468
rect 29052 72428 29058 72440
rect 237742 72428 237748 72440
rect 237800 72428 237806 72480
rect 328822 72428 328828 72480
rect 328880 72468 328886 72480
rect 470594 72468 470600 72480
rect 328880 72440 470600 72468
rect 328880 72428 328886 72440
rect 470594 72428 470600 72440
rect 470652 72428 470658 72480
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 230014 71720 230020 71732
rect 3384 71692 230020 71720
rect 3384 71680 3390 71692
rect 230014 71680 230020 71692
rect 230072 71680 230078 71732
rect 310606 71136 310612 71188
rect 310664 71176 310670 71188
rect 382274 71176 382280 71188
rect 310664 71148 382280 71176
rect 310664 71136 310670 71148
rect 382274 71136 382280 71148
rect 382332 71136 382338 71188
rect 201586 71068 201592 71120
rect 201644 71108 201650 71120
rect 273438 71108 273444 71120
rect 201644 71080 273444 71108
rect 201644 71068 201650 71080
rect 273438 71068 273444 71080
rect 273496 71068 273502 71120
rect 325878 71068 325884 71120
rect 325936 71108 325942 71120
rect 456886 71108 456892 71120
rect 325936 71080 456892 71108
rect 325936 71068 325942 71080
rect 456886 71068 456892 71080
rect 456944 71068 456950 71120
rect 121454 71000 121460 71052
rect 121512 71040 121518 71052
rect 257062 71040 257068 71052
rect 121512 71012 257068 71040
rect 121512 71000 121518 71012
rect 257062 71000 257068 71012
rect 257120 71000 257126 71052
rect 303798 71000 303804 71052
rect 303856 71040 303862 71052
rect 349154 71040 349160 71052
rect 303856 71012 349160 71040
rect 303856 71000 303862 71012
rect 349154 71000 349160 71012
rect 349212 71000 349218 71052
rect 349798 71000 349804 71052
rect 349856 71040 349862 71052
rect 571978 71040 571984 71052
rect 349856 71012 571984 71040
rect 349856 71000 349862 71012
rect 571978 71000 571984 71012
rect 572036 71000 572042 71052
rect 209866 69776 209872 69828
rect 209924 69816 209930 69828
rect 275094 69816 275100 69828
rect 209924 69788 275100 69816
rect 209924 69776 209930 69788
rect 275094 69776 275100 69788
rect 275152 69776 275158 69828
rect 309134 69776 309140 69828
rect 309192 69816 309198 69828
rect 374086 69816 374092 69828
rect 309192 69788 374092 69816
rect 309192 69776 309198 69788
rect 374086 69776 374092 69788
rect 374144 69776 374150 69828
rect 157334 69708 157340 69760
rect 157392 69748 157398 69760
rect 264330 69748 264336 69760
rect 157392 69720 264336 69748
rect 157392 69708 157398 69720
rect 264330 69708 264336 69720
rect 264388 69708 264394 69760
rect 321554 69708 321560 69760
rect 321612 69748 321618 69760
rect 434714 69748 434720 69760
rect 321612 69720 434720 69748
rect 321612 69708 321618 69720
rect 434714 69708 434720 69720
rect 434772 69708 434778 69760
rect 110414 69640 110420 69692
rect 110472 69680 110478 69692
rect 254762 69680 254768 69692
rect 110472 69652 254768 69680
rect 110472 69640 110478 69652
rect 254762 69640 254768 69652
rect 254820 69640 254826 69692
rect 302602 69640 302608 69692
rect 302660 69680 302666 69692
rect 342254 69680 342260 69692
rect 302660 69652 342260 69680
rect 302660 69640 302666 69652
rect 342254 69640 342260 69652
rect 342312 69640 342318 69692
rect 352650 69640 352656 69692
rect 352708 69680 352714 69692
rect 575474 69680 575480 69692
rect 352708 69652 575480 69680
rect 352708 69640 352714 69652
rect 575474 69640 575480 69652
rect 575532 69640 575538 69692
rect 216674 68416 216680 68468
rect 216732 68456 216738 68468
rect 276474 68456 276480 68468
rect 216732 68428 276480 68456
rect 216732 68416 216738 68428
rect 276474 68416 276480 68428
rect 276532 68416 276538 68468
rect 314746 68416 314752 68468
rect 314804 68456 314810 68468
rect 401594 68456 401600 68468
rect 314804 68428 401600 68456
rect 314804 68416 314810 68428
rect 401594 68416 401600 68428
rect 401652 68416 401658 68468
rect 161474 68348 161480 68400
rect 161532 68388 161538 68400
rect 265250 68388 265256 68400
rect 161532 68360 265256 68388
rect 161532 68348 161538 68360
rect 265250 68348 265256 68360
rect 265308 68348 265314 68400
rect 332042 68348 332048 68400
rect 332100 68388 332106 68400
rect 476114 68388 476120 68400
rect 332100 68360 476120 68388
rect 332100 68348 332106 68360
rect 476114 68348 476120 68360
rect 476172 68348 476178 68400
rect 93854 68280 93860 68332
rect 93912 68320 93918 68332
rect 251174 68320 251180 68332
rect 93912 68292 251180 68320
rect 93912 68280 93918 68292
rect 251174 68280 251180 68292
rect 251232 68280 251238 68332
rect 335630 68280 335636 68332
rect 335688 68320 335694 68332
rect 503714 68320 503720 68332
rect 335688 68292 503720 68320
rect 335688 68280 335694 68292
rect 503714 68280 503720 68292
rect 503772 68280 503778 68332
rect 165614 66988 165620 67040
rect 165672 67028 165678 67040
rect 266078 67028 266084 67040
rect 165672 67000 266084 67028
rect 165672 66988 165678 67000
rect 266078 66988 266084 67000
rect 266136 66988 266142 67040
rect 315390 66988 315396 67040
rect 315448 67028 315454 67040
rect 405734 67028 405740 67040
rect 315448 67000 405740 67028
rect 315448 66988 315454 67000
rect 405734 66988 405740 67000
rect 405792 66988 405798 67040
rect 95234 66920 95240 66972
rect 95292 66960 95298 66972
rect 251726 66960 251732 66972
rect 95292 66932 251732 66960
rect 95292 66920 95298 66932
rect 251726 66920 251732 66932
rect 251784 66920 251790 66972
rect 332594 66920 332600 66972
rect 332652 66960 332658 66972
rect 488534 66960 488540 66972
rect 332652 66932 488540 66960
rect 332652 66920 332658 66932
rect 488534 66920 488540 66932
rect 488592 66920 488598 66972
rect 69014 66852 69020 66904
rect 69072 66892 69078 66904
rect 246022 66892 246028 66904
rect 69072 66864 246028 66892
rect 69072 66852 69078 66864
rect 246022 66852 246028 66864
rect 246080 66852 246086 66904
rect 265066 66852 265072 66904
rect 265124 66892 265130 66904
rect 286502 66892 286508 66904
rect 265124 66864 286508 66892
rect 265124 66852 265130 66864
rect 286502 66852 286508 66864
rect 286560 66852 286566 66904
rect 296714 66852 296720 66904
rect 296772 66892 296778 66904
rect 314746 66892 314752 66904
rect 296772 66864 314752 66892
rect 296772 66852 296778 66864
rect 314746 66852 314752 66864
rect 314804 66852 314810 66904
rect 342346 66852 342352 66904
rect 342404 66892 342410 66904
rect 535454 66892 535460 66904
rect 342404 66864 535460 66892
rect 342404 66852 342410 66864
rect 535454 66852 535460 66864
rect 535512 66852 535518 66904
rect 172514 65628 172520 65680
rect 172572 65668 172578 65680
rect 267458 65668 267464 65680
rect 172572 65640 267464 65668
rect 172572 65628 172578 65640
rect 267458 65628 267464 65640
rect 267516 65628 267522 65680
rect 318334 65628 318340 65680
rect 318392 65668 318398 65680
rect 419534 65668 419540 65680
rect 318392 65640 419540 65668
rect 318392 65628 318398 65640
rect 419534 65628 419540 65640
rect 419592 65628 419598 65680
rect 82814 65560 82820 65612
rect 82872 65600 82878 65612
rect 248690 65600 248696 65612
rect 82872 65572 248696 65600
rect 82872 65560 82878 65572
rect 248690 65560 248696 65572
rect 248748 65560 248754 65612
rect 333974 65560 333980 65612
rect 334032 65600 334038 65612
rect 495434 65600 495440 65612
rect 334032 65572 495440 65600
rect 334032 65560 334038 65572
rect 495434 65560 495440 65572
rect 495492 65560 495498 65612
rect 44174 65492 44180 65544
rect 44232 65532 44238 65544
rect 241238 65532 241244 65544
rect 44232 65504 241244 65532
rect 44232 65492 44238 65504
rect 241238 65492 241244 65504
rect 241296 65492 241302 65544
rect 348050 65492 348056 65544
rect 348108 65532 348114 65544
rect 563698 65532 563704 65544
rect 348108 65504 563704 65532
rect 348108 65492 348114 65504
rect 563698 65492 563704 65504
rect 563756 65492 563762 65544
rect 179414 64268 179420 64320
rect 179472 64308 179478 64320
rect 270126 64308 270132 64320
rect 179472 64280 270132 64308
rect 179472 64268 179478 64280
rect 270126 64268 270132 64280
rect 270184 64268 270190 64320
rect 316034 64268 316040 64320
rect 316092 64308 316098 64320
rect 407114 64308 407120 64320
rect 316092 64280 407120 64308
rect 316092 64268 316098 64280
rect 407114 64268 407120 64280
rect 407172 64268 407178 64320
rect 88334 64200 88340 64252
rect 88392 64240 88398 64252
rect 250254 64240 250260 64252
rect 88392 64212 250260 64240
rect 88392 64200 88398 64212
rect 250254 64200 250260 64212
rect 250312 64200 250318 64252
rect 319530 64200 319536 64252
rect 319588 64240 319594 64252
rect 426434 64240 426440 64252
rect 319588 64212 426440 64240
rect 319588 64200 319594 64212
rect 426434 64200 426440 64212
rect 426492 64200 426498 64252
rect 57974 64132 57980 64184
rect 58032 64172 58038 64184
rect 243814 64172 243820 64184
rect 58032 64144 243820 64172
rect 58032 64132 58038 64144
rect 243814 64132 243820 64144
rect 243872 64132 243878 64184
rect 341242 64132 341248 64184
rect 341300 64172 341306 64184
rect 531314 64172 531320 64184
rect 341300 64144 531320 64172
rect 341300 64132 341306 64144
rect 531314 64132 531320 64144
rect 531372 64132 531378 64184
rect 183554 62908 183560 62960
rect 183612 62948 183618 62960
rect 269666 62948 269672 62960
rect 183612 62920 269672 62948
rect 183612 62908 183618 62920
rect 269666 62908 269672 62920
rect 269724 62908 269730 62960
rect 307846 62908 307852 62960
rect 307904 62948 307910 62960
rect 372614 62948 372620 62960
rect 307904 62920 372620 62948
rect 307904 62908 307910 62920
rect 372614 62908 372620 62920
rect 372672 62908 372678 62960
rect 74534 62840 74540 62892
rect 74592 62880 74598 62892
rect 247402 62880 247408 62892
rect 74592 62852 247408 62880
rect 74592 62840 74598 62852
rect 247402 62840 247408 62852
rect 247460 62840 247466 62892
rect 321002 62840 321008 62892
rect 321060 62880 321066 62892
rect 433334 62880 433340 62892
rect 321060 62852 433340 62880
rect 321060 62840 321066 62852
rect 433334 62840 433340 62852
rect 433392 62840 433398 62892
rect 64874 62772 64880 62824
rect 64932 62812 64938 62824
rect 242158 62812 242164 62824
rect 64932 62784 242164 62812
rect 64932 62772 64938 62784
rect 242158 62772 242164 62784
rect 242216 62772 242222 62824
rect 345566 62772 345572 62824
rect 345624 62812 345630 62824
rect 552014 62812 552020 62824
rect 345624 62784 552020 62812
rect 345624 62772 345630 62784
rect 552014 62772 552020 62784
rect 552072 62772 552078 62824
rect 186314 61480 186320 61532
rect 186372 61520 186378 61532
rect 271322 61520 271328 61532
rect 186372 61492 271328 61520
rect 186372 61480 186378 61492
rect 271322 61480 271328 61492
rect 271380 61480 271386 61532
rect 306466 61480 306472 61532
rect 306524 61520 306530 61532
rect 361574 61520 361580 61532
rect 306524 61492 361580 61520
rect 306524 61480 306530 61492
rect 361574 61480 361580 61492
rect 361632 61480 361638 61532
rect 63494 61412 63500 61464
rect 63552 61452 63558 61464
rect 245102 61452 245108 61464
rect 63552 61424 245108 61452
rect 63552 61412 63558 61424
rect 245102 61412 245108 61424
rect 245160 61412 245166 61464
rect 335998 61412 336004 61464
rect 336056 61452 336062 61464
rect 437474 61452 437480 61464
rect 336056 61424 437480 61452
rect 336056 61412 336062 61424
rect 437474 61412 437480 61424
rect 437532 61412 437538 61464
rect 11054 61344 11060 61396
rect 11112 61384 11118 61396
rect 232498 61384 232504 61396
rect 11112 61356 232504 61384
rect 11112 61344 11118 61356
rect 232498 61344 232504 61356
rect 232556 61344 232562 61396
rect 346394 61344 346400 61396
rect 346452 61384 346458 61396
rect 556154 61384 556160 61396
rect 346452 61356 556160 61384
rect 346452 61344 346458 61356
rect 556154 61344 556160 61356
rect 556212 61344 556218 61396
rect 354306 60664 354312 60716
rect 354364 60704 354370 60716
rect 580166 60704 580172 60716
rect 354364 60676 580172 60704
rect 354364 60664 354370 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 208394 60120 208400 60172
rect 208452 60160 208458 60172
rect 273990 60160 273996 60172
rect 208452 60132 273996 60160
rect 208452 60120 208458 60132
rect 273990 60120 273996 60132
rect 274048 60120 274054 60172
rect 301130 60120 301136 60172
rect 301188 60160 301194 60172
rect 335446 60160 335452 60172
rect 301188 60132 335452 60160
rect 301188 60120 301194 60132
rect 335446 60120 335452 60132
rect 335504 60120 335510 60172
rect 149054 60052 149060 60104
rect 149112 60092 149118 60104
rect 262674 60092 262680 60104
rect 149112 60064 262680 60092
rect 149112 60052 149118 60064
rect 262674 60052 262680 60064
rect 262732 60052 262738 60104
rect 313550 60052 313556 60104
rect 313608 60092 313614 60104
rect 396074 60092 396080 60104
rect 313608 60064 396080 60092
rect 313608 60052 313614 60064
rect 396074 60052 396080 60064
rect 396132 60052 396138 60104
rect 12434 59984 12440 60036
rect 12492 60024 12498 60036
rect 234798 60024 234804 60036
rect 12492 59996 234804 60024
rect 12492 59984 12498 59996
rect 234798 59984 234804 59996
rect 234856 59984 234862 60036
rect 318886 59984 318892 60036
rect 318944 60024 318950 60036
rect 422294 60024 422300 60036
rect 318944 59996 422300 60024
rect 318944 59984 318950 59996
rect 422294 59984 422300 59996
rect 422352 59984 422358 60036
rect 222194 58760 222200 58812
rect 222252 58800 222258 58812
rect 277762 58800 277768 58812
rect 222252 58772 277768 58800
rect 222252 58760 222258 58772
rect 277762 58760 277768 58772
rect 277820 58760 277826 58812
rect 321830 58760 321836 58812
rect 321888 58800 321894 58812
rect 436094 58800 436100 58812
rect 321888 58772 436100 58800
rect 321888 58760 321894 58772
rect 436094 58760 436100 58772
rect 436152 58760 436158 58812
rect 131114 58692 131120 58744
rect 131172 58732 131178 58744
rect 258994 58732 259000 58744
rect 131172 58704 259000 58732
rect 131172 58692 131178 58704
rect 258994 58692 259000 58704
rect 259052 58692 259058 58744
rect 323486 58692 323492 58744
rect 323544 58732 323550 58744
rect 444374 58732 444380 58744
rect 323544 58704 444380 58732
rect 323544 58692 323550 58704
rect 444374 58692 444380 58704
rect 444432 58692 444438 58744
rect 84194 58624 84200 58676
rect 84252 58664 84258 58676
rect 249242 58664 249248 58676
rect 84252 58636 249248 58664
rect 84252 58624 84258 58636
rect 249242 58624 249248 58636
rect 249300 58624 249306 58676
rect 298462 58624 298468 58676
rect 298520 58664 298526 58676
rect 323026 58664 323032 58676
rect 298520 58636 323032 58664
rect 298520 58624 298526 58636
rect 323026 58624 323032 58636
rect 323084 58624 323090 58676
rect 349246 58624 349252 58676
rect 349304 58664 349310 58676
rect 569954 58664 569960 58676
rect 349304 58636 569960 58664
rect 349304 58624 349310 58636
rect 569954 58624 569960 58636
rect 570012 58624 570018 58676
rect 314930 57332 314936 57384
rect 314988 57372 314994 57384
rect 402974 57372 402980 57384
rect 314988 57344 402980 57372
rect 314988 57332 314994 57344
rect 402974 57332 402980 57344
rect 403032 57332 403038 57384
rect 133874 57264 133880 57316
rect 133932 57304 133938 57316
rect 259638 57304 259644 57316
rect 133932 57276 259644 57304
rect 133932 57264 133938 57276
rect 259638 57264 259644 57276
rect 259696 57264 259702 57316
rect 324866 57264 324872 57316
rect 324924 57304 324930 57316
rect 451274 57304 451280 57316
rect 324924 57276 451280 57304
rect 324924 57264 324930 57276
rect 451274 57264 451280 57276
rect 451332 57264 451338 57316
rect 73154 57196 73160 57248
rect 73212 57236 73218 57248
rect 247034 57236 247040 57248
rect 73212 57208 247040 57236
rect 73212 57196 73218 57208
rect 247034 57196 247040 57208
rect 247092 57196 247098 57248
rect 338574 57196 338580 57248
rect 338632 57236 338638 57248
rect 517514 57236 517520 57248
rect 338632 57208 517520 57236
rect 338632 57196 338638 57208
rect 517514 57196 517520 57208
rect 517572 57196 517578 57248
rect 317874 55972 317880 56024
rect 317932 56012 317938 56024
rect 416774 56012 416780 56024
rect 317932 55984 416780 56012
rect 317932 55972 317938 55984
rect 416774 55972 416780 55984
rect 416832 55972 416838 56024
rect 143626 55904 143632 55956
rect 143684 55944 143690 55956
rect 261662 55944 261668 55956
rect 143684 55916 261668 55944
rect 143684 55904 143690 55916
rect 261662 55904 261668 55916
rect 261720 55904 261726 55956
rect 327166 55904 327172 55956
rect 327224 55944 327230 55956
rect 462314 55944 462320 55956
rect 327224 55916 462320 55944
rect 327224 55904 327230 55916
rect 462314 55904 462320 55916
rect 462372 55904 462378 55956
rect 62114 55836 62120 55888
rect 62172 55876 62178 55888
rect 244826 55876 244832 55888
rect 62172 55848 244832 55876
rect 62172 55836 62178 55848
rect 244826 55836 244832 55848
rect 244884 55836 244890 55888
rect 343726 55836 343732 55888
rect 343784 55876 343790 55888
rect 542354 55876 542360 55888
rect 343784 55848 542360 55876
rect 343784 55836 343790 55848
rect 542354 55836 542360 55848
rect 542412 55836 542418 55888
rect 320174 54612 320180 54664
rect 320232 54652 320238 54664
rect 427814 54652 427820 54664
rect 320232 54624 427820 54652
rect 320232 54612 320238 54624
rect 427814 54612 427820 54624
rect 427872 54612 427878 54664
rect 127066 54544 127072 54596
rect 127124 54584 127130 54596
rect 258442 54584 258448 54596
rect 127124 54556 258448 54584
rect 127124 54544 127130 54556
rect 258442 54544 258448 54556
rect 258500 54544 258506 54596
rect 327810 54544 327816 54596
rect 327868 54584 327874 54596
rect 465166 54584 465172 54596
rect 327868 54556 465172 54584
rect 327868 54544 327874 54556
rect 465166 54544 465172 54556
rect 465224 54544 465230 54596
rect 77294 54476 77300 54528
rect 77352 54516 77358 54528
rect 247218 54516 247224 54528
rect 77352 54488 247224 54516
rect 77352 54476 77358 54488
rect 247218 54476 247224 54488
rect 247276 54476 247282 54528
rect 349706 54476 349712 54528
rect 349764 54516 349770 54528
rect 574094 54516 574100 54528
rect 349764 54488 574100 54516
rect 349764 54476 349770 54488
rect 574094 54476 574100 54488
rect 574152 54476 574158 54528
rect 162854 53116 162860 53168
rect 162912 53156 162918 53168
rect 265158 53156 265164 53168
rect 162912 53128 265164 53156
rect 162912 53116 162918 53128
rect 265158 53116 265164 53128
rect 265216 53116 265222 53168
rect 324498 53116 324504 53168
rect 324556 53156 324562 53168
rect 448606 53156 448612 53168
rect 324556 53128 448612 53156
rect 324556 53116 324562 53128
rect 448606 53116 448612 53128
rect 448664 53116 448670 53168
rect 114554 53048 114560 53100
rect 114612 53088 114618 53100
rect 255590 53088 255596 53100
rect 114612 53060 255596 53088
rect 114612 53048 114618 53060
rect 255590 53048 255596 53060
rect 255648 53048 255654 53100
rect 300302 53048 300308 53100
rect 300360 53088 300366 53100
rect 332594 53088 332600 53100
rect 300360 53060 332600 53088
rect 300360 53048 300366 53060
rect 332594 53048 332600 53060
rect 332652 53048 332658 53100
rect 333238 53048 333244 53100
rect 333296 53088 333302 53100
rect 469214 53088 469220 53100
rect 333296 53060 469220 53088
rect 333296 53048 333302 53060
rect 469214 53048 469220 53060
rect 469272 53048 469278 53100
rect 166994 51756 167000 51808
rect 167052 51796 167058 51808
rect 266446 51796 266452 51808
rect 167052 51768 266452 51796
rect 167052 51756 167058 51768
rect 266446 51756 266452 51768
rect 266504 51756 266510 51808
rect 322198 51756 322204 51808
rect 322256 51796 322262 51808
rect 438854 51796 438860 51808
rect 322256 51768 438860 51796
rect 322256 51756 322262 51768
rect 438854 51756 438860 51768
rect 438912 51756 438918 51808
rect 8294 51688 8300 51740
rect 8352 51728 8358 51740
rect 233694 51728 233700 51740
rect 8352 51700 233700 51728
rect 8352 51688 8358 51700
rect 233694 51688 233700 51700
rect 233752 51688 233758 51740
rect 329282 51688 329288 51740
rect 329340 51728 329346 51740
rect 473354 51728 473360 51740
rect 329340 51700 473360 51728
rect 329340 51688 329346 51700
rect 473354 51688 473360 51700
rect 473412 51688 473418 51740
rect 169754 50396 169760 50448
rect 169812 50436 169818 50448
rect 266722 50436 266728 50448
rect 169812 50408 266728 50436
rect 169812 50396 169818 50408
rect 266722 50396 266728 50408
rect 266780 50396 266786 50448
rect 323670 50396 323676 50448
rect 323728 50436 323734 50448
rect 445754 50436 445760 50448
rect 323728 50408 445760 50436
rect 323728 50396 323734 50408
rect 445754 50396 445760 50408
rect 445812 50396 445818 50448
rect 66254 50328 66260 50380
rect 66312 50368 66318 50380
rect 245746 50368 245752 50380
rect 66312 50340 245752 50368
rect 66312 50328 66318 50340
rect 245746 50328 245752 50340
rect 245804 50328 245810 50380
rect 331674 50328 331680 50380
rect 331732 50368 331738 50380
rect 484394 50368 484400 50380
rect 331732 50340 484400 50368
rect 331732 50328 331738 50340
rect 484394 50328 484400 50340
rect 484452 50328 484458 50380
rect 229094 49104 229100 49156
rect 229152 49144 229158 49156
rect 275370 49144 275376 49156
rect 229152 49116 275376 49144
rect 229152 49104 229158 49116
rect 275370 49104 275376 49116
rect 275428 49104 275434 49156
rect 111794 49036 111800 49088
rect 111852 49076 111858 49088
rect 255038 49076 255044 49088
rect 111852 49048 255044 49076
rect 111852 49036 111858 49048
rect 255038 49036 255044 49048
rect 255096 49036 255102 49088
rect 331306 49036 331312 49088
rect 331364 49076 331370 49088
rect 481726 49076 481732 49088
rect 331364 49048 481732 49076
rect 331364 49036 331370 49048
rect 481726 49036 481732 49048
rect 481784 49036 481790 49088
rect 2774 48968 2780 49020
rect 2832 49008 2838 49020
rect 232590 49008 232596 49020
rect 2832 48980 232596 49008
rect 2832 48968 2838 48980
rect 232590 48968 232596 48980
rect 232648 48968 232654 49020
rect 333146 48968 333152 49020
rect 333204 49008 333210 49020
rect 491294 49008 491300 49020
rect 333204 48980 491300 49008
rect 333204 48968 333210 48980
rect 491294 48968 491300 48980
rect 491352 48968 491358 49020
rect 176654 47608 176660 47660
rect 176712 47648 176718 47660
rect 267918 47648 267924 47660
rect 176712 47620 267924 47648
rect 176712 47608 176718 47620
rect 267918 47608 267924 47620
rect 267976 47608 267982 47660
rect 334618 47608 334624 47660
rect 334676 47648 334682 47660
rect 498286 47648 498292 47660
rect 334676 47620 498292 47648
rect 334676 47608 334682 47620
rect 498286 47608 498292 47620
rect 498344 47608 498350 47660
rect 59354 47540 59360 47592
rect 59412 47580 59418 47592
rect 243538 47580 243544 47592
rect 59412 47552 243544 47580
rect 59412 47540 59418 47552
rect 243538 47540 243544 47552
rect 243596 47540 243602 47592
rect 337102 47540 337108 47592
rect 337160 47580 337166 47592
rect 510614 47580 510620 47592
rect 337160 47552 510620 47580
rect 337160 47540 337166 47552
rect 510614 47540 510620 47552
rect 510672 47540 510678 47592
rect 354214 46860 354220 46912
rect 354272 46900 354278 46912
rect 580166 46900 580172 46912
rect 354272 46872 580172 46900
rect 354272 46860 354278 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 187694 46316 187700 46368
rect 187752 46356 187758 46368
rect 270678 46356 270684 46368
rect 187752 46328 270684 46356
rect 187752 46316 187758 46328
rect 270678 46316 270684 46328
rect 270736 46316 270742 46368
rect 99374 46248 99380 46300
rect 99432 46288 99438 46300
rect 252830 46288 252836 46300
rect 99432 46260 252836 46288
rect 99432 46248 99438 46260
rect 252830 46248 252836 46260
rect 252888 46248 252894 46300
rect 303982 46248 303988 46300
rect 304040 46288 304046 46300
rect 349246 46288 349252 46300
rect 304040 46260 349252 46288
rect 304040 46248 304046 46260
rect 349246 46248 349252 46260
rect 349304 46248 349310 46300
rect 33134 46180 33140 46232
rect 33192 46220 33198 46232
rect 238846 46220 238852 46232
rect 33192 46192 238852 46220
rect 33192 46180 33198 46192
rect 238846 46180 238852 46192
rect 238904 46180 238910 46232
rect 334342 46180 334348 46232
rect 334400 46220 334406 46232
rect 499574 46220 499580 46232
rect 334400 46192 499580 46220
rect 334400 46180 334406 46192
rect 499574 46180 499580 46192
rect 499632 46180 499638 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 229922 45540 229928 45552
rect 3568 45512 229928 45540
rect 3568 45500 3574 45512
rect 229922 45500 229928 45512
rect 229980 45500 229986 45552
rect 226334 44888 226340 44940
rect 226392 44928 226398 44940
rect 278866 44928 278872 44940
rect 226392 44900 278872 44928
rect 226392 44888 226398 44900
rect 278866 44888 278872 44900
rect 278924 44888 278930 44940
rect 335538 44888 335544 44940
rect 335596 44928 335602 44940
rect 502334 44928 502340 44940
rect 335596 44900 502340 44928
rect 335596 44888 335602 44900
rect 502334 44888 502340 44900
rect 502392 44888 502398 44940
rect 60826 44820 60832 44872
rect 60884 44860 60890 44872
rect 244550 44860 244556 44872
rect 60884 44832 244556 44860
rect 60884 44820 60890 44832
rect 244550 44820 244556 44832
rect 244608 44820 244614 44872
rect 338758 44820 338764 44872
rect 338816 44860 338822 44872
rect 521654 44860 521660 44872
rect 338816 44832 521660 44860
rect 338816 44820 338822 44832
rect 521654 44820 521660 44832
rect 521712 44820 521718 44872
rect 191834 43460 191840 43512
rect 191892 43500 191898 43512
rect 270586 43500 270592 43512
rect 191892 43472 270592 43500
rect 191892 43460 191898 43472
rect 270586 43460 270592 43472
rect 270644 43460 270650 43512
rect 335814 43460 335820 43512
rect 335872 43500 335878 43512
rect 506474 43500 506480 43512
rect 335872 43472 506480 43500
rect 335872 43460 335878 43472
rect 506474 43460 506480 43472
rect 506532 43460 506538 43512
rect 48314 43392 48320 43444
rect 48372 43432 48378 43444
rect 241974 43432 241980 43444
rect 48372 43404 241980 43432
rect 48372 43392 48378 43404
rect 241974 43392 241980 43404
rect 242032 43392 242038 43444
rect 340046 43392 340052 43444
rect 340104 43432 340110 43444
rect 524414 43432 524420 43444
rect 340104 43404 524420 43432
rect 340104 43392 340110 43404
rect 524414 43392 524420 43404
rect 524472 43392 524478 43444
rect 194594 42168 194600 42220
rect 194652 42208 194658 42220
rect 272150 42208 272156 42220
rect 194652 42180 272156 42208
rect 194652 42168 194658 42180
rect 272150 42168 272156 42180
rect 272208 42168 272214 42220
rect 110506 42100 110512 42152
rect 110564 42140 110570 42152
rect 254578 42140 254584 42152
rect 110564 42112 254584 42140
rect 110564 42100 110570 42112
rect 254578 42100 254584 42112
rect 254636 42100 254642 42152
rect 336918 42100 336924 42152
rect 336976 42140 336982 42152
rect 509234 42140 509240 42152
rect 336976 42112 509240 42140
rect 336976 42100 336982 42112
rect 509234 42100 509240 42112
rect 509292 42100 509298 42152
rect 52454 42032 52460 42084
rect 52512 42072 52518 42084
rect 242618 42072 242624 42084
rect 52512 42044 242624 42072
rect 52512 42032 52518 42044
rect 242618 42032 242624 42044
rect 242676 42032 242682 42084
rect 301314 42032 301320 42084
rect 301372 42072 301378 42084
rect 336734 42072 336740 42084
rect 301372 42044 336740 42072
rect 301372 42032 301378 42044
rect 336734 42032 336740 42044
rect 336792 42032 336798 42084
rect 341886 42032 341892 42084
rect 341944 42072 341950 42084
rect 528554 42072 528560 42084
rect 341944 42044 528560 42072
rect 341944 42032 341950 42044
rect 528554 42032 528560 42044
rect 528612 42032 528618 42084
rect 205634 40808 205640 40860
rect 205692 40848 205698 40860
rect 274266 40848 274272 40860
rect 205692 40820 274272 40848
rect 205692 40808 205698 40820
rect 274266 40808 274272 40820
rect 274324 40808 274330 40860
rect 81434 40740 81440 40792
rect 81492 40780 81498 40792
rect 248782 40780 248788 40792
rect 81492 40752 248788 40780
rect 81492 40740 81498 40752
rect 248782 40740 248788 40752
rect 248840 40740 248846 40792
rect 337286 40740 337292 40792
rect 337344 40780 337350 40792
rect 513374 40780 513380 40792
rect 337344 40752 513380 40780
rect 337344 40740 337350 40752
rect 513374 40740 513380 40752
rect 513432 40740 513438 40792
rect 44266 40672 44272 40724
rect 44324 40712 44330 40724
rect 224310 40712 224316 40724
rect 44324 40684 224316 40712
rect 44324 40672 44330 40684
rect 224310 40672 224316 40684
rect 224368 40672 224374 40724
rect 342898 40672 342904 40724
rect 342956 40712 342962 40724
rect 539686 40712 539692 40724
rect 342956 40684 539692 40712
rect 342956 40672 342962 40684
rect 539686 40672 539692 40684
rect 539744 40672 539750 40724
rect 223574 39448 223580 39500
rect 223632 39488 223638 39500
rect 276658 39488 276664 39500
rect 223632 39460 276664 39488
rect 223632 39448 223638 39460
rect 276658 39448 276664 39460
rect 276716 39448 276722 39500
rect 302786 39448 302792 39500
rect 302844 39488 302850 39500
rect 343726 39488 343732 39500
rect 302844 39460 343732 39488
rect 302844 39448 302850 39460
rect 343726 39448 343732 39460
rect 343784 39448 343790 39500
rect 67634 39380 67640 39432
rect 67692 39420 67698 39432
rect 245838 39420 245844 39432
rect 67692 39392 245844 39420
rect 67692 39380 67698 39392
rect 245838 39380 245844 39392
rect 245896 39380 245902 39432
rect 338298 39380 338304 39432
rect 338356 39420 338362 39432
rect 516134 39420 516140 39432
rect 338356 39392 516140 39420
rect 338356 39380 338362 39392
rect 516134 39380 516140 39392
rect 516192 39380 516198 39432
rect 6914 39312 6920 39364
rect 6972 39352 6978 39364
rect 231118 39352 231124 39364
rect 6972 39324 231124 39352
rect 6972 39312 6978 39324
rect 231118 39312 231124 39324
rect 231176 39312 231182 39364
rect 343634 39312 343640 39364
rect 343692 39352 343698 39364
rect 546494 39352 546500 39364
rect 343692 39324 546500 39352
rect 343692 39312 343698 39324
rect 546494 39312 546500 39324
rect 546552 39312 546558 39364
rect 135346 37952 135352 38004
rect 135404 37992 135410 38004
rect 259822 37992 259828 38004
rect 135404 37964 259828 37992
rect 135404 37952 135410 37964
rect 259822 37952 259828 37964
rect 259880 37952 259886 38004
rect 338482 37952 338488 38004
rect 338540 37992 338546 38004
rect 520274 37992 520280 38004
rect 338540 37964 520280 37992
rect 338540 37952 338546 37964
rect 520274 37952 520280 37964
rect 520332 37952 520338 38004
rect 102134 37884 102140 37936
rect 102192 37924 102198 37936
rect 253014 37924 253020 37936
rect 102192 37896 253020 37924
rect 102192 37884 102198 37896
rect 253014 37884 253020 37896
rect 253072 37884 253078 37936
rect 345106 37884 345112 37936
rect 345164 37924 345170 37936
rect 549254 37924 549260 37936
rect 345164 37896 549260 37924
rect 345164 37884 345170 37896
rect 549254 37884 549260 37896
rect 549312 37884 549318 37936
rect 138014 36592 138020 36644
rect 138072 36632 138078 36644
rect 259914 36632 259920 36644
rect 138072 36604 259920 36632
rect 138072 36592 138078 36604
rect 259914 36592 259920 36604
rect 259972 36592 259978 36644
rect 339954 36592 339960 36644
rect 340012 36632 340018 36644
rect 527174 36632 527180 36644
rect 340012 36604 527180 36632
rect 340012 36592 340018 36604
rect 527174 36592 527180 36604
rect 527232 36592 527238 36644
rect 22094 36524 22100 36576
rect 22152 36564 22158 36576
rect 235258 36564 235264 36576
rect 22152 36536 235264 36564
rect 22152 36524 22158 36536
rect 235258 36524 235264 36536
rect 235316 36524 235322 36576
rect 345290 36524 345296 36576
rect 345348 36564 345354 36576
rect 553394 36564 553400 36576
rect 345348 36536 553400 36564
rect 345348 36524 345354 36536
rect 553394 36524 553400 36536
rect 553452 36524 553458 36576
rect 142154 35232 142160 35284
rect 142212 35272 142218 35284
rect 261202 35272 261208 35284
rect 142212 35244 261208 35272
rect 142212 35232 142218 35244
rect 261202 35232 261208 35244
rect 261260 35232 261266 35284
rect 341426 35232 341432 35284
rect 341484 35272 341490 35284
rect 534074 35272 534080 35284
rect 341484 35244 534080 35272
rect 341484 35232 341490 35244
rect 534074 35232 534080 35244
rect 534132 35232 534138 35284
rect 17954 35164 17960 35216
rect 18012 35204 18018 35216
rect 235350 35204 235356 35216
rect 18012 35176 235356 35204
rect 18012 35164 18018 35176
rect 235350 35164 235356 35176
rect 235408 35164 235414 35216
rect 346578 35164 346584 35216
rect 346636 35204 346642 35216
rect 556246 35204 556252 35216
rect 346636 35176 556252 35204
rect 346636 35164 346642 35176
rect 556246 35164 556252 35176
rect 556304 35164 556310 35216
rect 151906 33804 151912 33856
rect 151964 33844 151970 33856
rect 262582 33844 262588 33856
rect 151964 33816 262588 33844
rect 151964 33804 151970 33816
rect 262582 33804 262588 33816
rect 262640 33804 262646 33856
rect 342714 33804 342720 33856
rect 342772 33844 342778 33856
rect 538214 33844 538220 33856
rect 342772 33816 538220 33844
rect 342772 33804 342778 33816
rect 538214 33804 538220 33816
rect 538272 33804 538278 33856
rect 97994 33736 98000 33788
rect 98052 33776 98058 33788
rect 251358 33776 251364 33788
rect 98052 33748 251364 33776
rect 98052 33736 98058 33748
rect 251358 33736 251364 33748
rect 251416 33736 251422 33788
rect 348234 33736 348240 33788
rect 348292 33776 348298 33788
rect 567194 33776 567200 33788
rect 348292 33748 567200 33776
rect 348292 33736 348298 33748
rect 567194 33736 567200 33748
rect 567252 33736 567258 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 229830 33096 229836 33108
rect 3568 33068 229836 33096
rect 3568 33056 3574 33068
rect 229830 33056 229836 33068
rect 229888 33056 229894 33108
rect 354122 33056 354128 33108
rect 354180 33096 354186 33108
rect 580166 33096 580172 33108
rect 354180 33068 580172 33096
rect 354180 33056 354186 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 304166 32444 304172 32496
rect 304224 32484 304230 32496
rect 353294 32484 353300 32496
rect 304224 32456 353300 32484
rect 304224 32444 304230 32456
rect 353294 32444 353300 32456
rect 353352 32444 353358 32496
rect 118694 32376 118700 32428
rect 118752 32416 118758 32428
rect 256970 32416 256976 32428
rect 118752 32388 256976 32416
rect 118752 32376 118758 32388
rect 256970 32376 256976 32388
rect 257028 32376 257034 32428
rect 314194 32376 314200 32428
rect 314252 32416 314258 32428
rect 400214 32416 400220 32428
rect 314252 32388 400220 32416
rect 314252 32376 314258 32388
rect 400214 32376 400220 32388
rect 400272 32376 400278 32428
rect 304994 31152 305000 31204
rect 305052 31192 305058 31204
rect 354674 31192 354680 31204
rect 305052 31164 354680 31192
rect 305052 31152 305058 31164
rect 354674 31152 354680 31164
rect 354732 31152 354738 31204
rect 155954 31084 155960 31136
rect 156012 31124 156018 31136
rect 263778 31124 263784 31136
rect 156012 31096 263784 31124
rect 156012 31084 156018 31096
rect 263778 31084 263784 31096
rect 263836 31084 263842 31136
rect 318058 31084 318064 31136
rect 318116 31124 318122 31136
rect 418154 31124 418160 31136
rect 318116 31096 418160 31124
rect 318116 31084 318122 31096
rect 418154 31084 418160 31096
rect 418212 31084 418218 31136
rect 109034 31016 109040 31068
rect 109092 31056 109098 31068
rect 254394 31056 254400 31068
rect 109092 31028 254400 31056
rect 109092 31016 109098 31028
rect 254394 31016 254400 31028
rect 254452 31016 254458 31068
rect 342622 31016 342628 31068
rect 342680 31056 342686 31068
rect 540974 31056 540980 31068
rect 342680 31028 540980 31056
rect 342680 31016 342686 31028
rect 540974 31016 540980 31028
rect 541032 31016 541038 31068
rect 160186 29656 160192 29708
rect 160244 29696 160250 29708
rect 264974 29696 264980 29708
rect 160244 29668 264980 29696
rect 160244 29656 160250 29668
rect 264974 29656 264980 29668
rect 265032 29656 265038 29708
rect 315114 29656 315120 29708
rect 315172 29696 315178 29708
rect 404354 29696 404360 29708
rect 315172 29668 404360 29696
rect 315172 29656 315178 29668
rect 404354 29656 404360 29668
rect 404412 29656 404418 29708
rect 104894 29588 104900 29640
rect 104952 29628 104958 29640
rect 253566 29628 253572 29640
rect 104952 29600 253572 29628
rect 104952 29588 104958 29600
rect 253566 29588 253572 29600
rect 253624 29588 253630 29640
rect 301774 29588 301780 29640
rect 301832 29628 301838 29640
rect 340966 29628 340972 29640
rect 301832 29600 340972 29628
rect 301832 29588 301838 29600
rect 340966 29588 340972 29600
rect 341024 29588 341030 29640
rect 345014 29588 345020 29640
rect 345072 29628 345078 29640
rect 547966 29628 547972 29640
rect 345072 29600 547972 29628
rect 345072 29588 345078 29600
rect 547966 29588 547972 29600
rect 548024 29588 548030 29640
rect 96614 28296 96620 28348
rect 96672 28336 96678 28348
rect 251910 28336 251916 28348
rect 96672 28308 251916 28336
rect 96672 28296 96678 28308
rect 251910 28296 251916 28308
rect 251968 28296 251974 28348
rect 316126 28296 316132 28348
rect 316184 28336 316190 28348
rect 411254 28336 411260 28348
rect 316184 28308 411260 28336
rect 316184 28296 316190 28308
rect 411254 28296 411260 28308
rect 411312 28296 411318 28348
rect 56594 28228 56600 28280
rect 56652 28268 56658 28280
rect 243354 28268 243360 28280
rect 56652 28240 243360 28268
rect 56652 28228 56658 28240
rect 243354 28228 243360 28240
rect 243412 28228 243418 28280
rect 302970 28228 302976 28280
rect 303028 28268 303034 28280
rect 346394 28268 346400 28280
rect 303028 28240 346400 28268
rect 303028 28228 303034 28240
rect 346394 28228 346400 28240
rect 346452 28228 346458 28280
rect 347038 28228 347044 28280
rect 347096 28268 347102 28280
rect 558914 28268 558920 28280
rect 347096 28240 558920 28268
rect 347096 28228 347102 28240
rect 558914 28228 558920 28240
rect 558972 28228 558978 28280
rect 212534 27004 212540 27056
rect 212592 27044 212598 27056
rect 275002 27044 275008 27056
rect 212592 27016 275008 27044
rect 212592 27004 212598 27016
rect 275002 27004 275008 27016
rect 275060 27004 275066 27056
rect 102226 26936 102232 26988
rect 102284 26976 102290 26988
rect 253106 26976 253112 26988
rect 102284 26948 253112 26976
rect 102284 26936 102290 26948
rect 253106 26936 253112 26948
rect 253164 26936 253170 26988
rect 310514 26936 310520 26988
rect 310572 26976 310578 26988
rect 382366 26976 382372 26988
rect 310572 26948 382372 26976
rect 310572 26936 310578 26948
rect 382366 26936 382372 26948
rect 382424 26936 382430 26988
rect 55214 26868 55220 26920
rect 55272 26908 55278 26920
rect 243446 26908 243452 26920
rect 55272 26880 243452 26908
rect 55272 26868 55278 26880
rect 243446 26868 243452 26880
rect 243504 26868 243510 26920
rect 300026 26868 300032 26920
rect 300084 26908 300090 26920
rect 332870 26908 332876 26920
rect 300084 26880 332876 26908
rect 300084 26868 300090 26880
rect 332870 26868 332876 26880
rect 332928 26868 332934 26920
rect 349430 26868 349436 26920
rect 349488 26908 349494 26920
rect 572806 26908 572812 26920
rect 349488 26880 572812 26908
rect 349488 26868 349494 26880
rect 572806 26868 572812 26880
rect 572864 26868 572870 26920
rect 185026 25576 185032 25628
rect 185084 25616 185090 25628
rect 269850 25616 269856 25628
rect 185084 25588 269856 25616
rect 185084 25576 185090 25588
rect 269850 25576 269856 25588
rect 269908 25576 269914 25628
rect 313918 25576 313924 25628
rect 313976 25616 313982 25628
rect 398926 25616 398932 25628
rect 313976 25588 398932 25616
rect 313976 25576 313982 25588
rect 398926 25576 398932 25588
rect 398984 25576 398990 25628
rect 86954 25508 86960 25560
rect 87012 25548 87018 25560
rect 249978 25548 249984 25560
rect 87012 25520 249984 25548
rect 87012 25508 87018 25520
rect 249978 25508 249984 25520
rect 250036 25508 250042 25560
rect 327350 25508 327356 25560
rect 327408 25548 327414 25560
rect 463694 25548 463700 25560
rect 327408 25520 463700 25548
rect 327408 25508 327414 25520
rect 463694 25508 463700 25520
rect 463752 25508 463758 25560
rect 154574 24148 154580 24200
rect 154632 24188 154638 24200
rect 264514 24188 264520 24200
rect 154632 24160 264520 24188
rect 154632 24148 154638 24160
rect 264514 24148 264520 24160
rect 264572 24148 264578 24200
rect 314654 24148 314660 24200
rect 314712 24188 314718 24200
rect 407206 24188 407212 24200
rect 314712 24160 407212 24188
rect 314712 24148 314718 24160
rect 407206 24148 407212 24160
rect 407264 24148 407270 24200
rect 27614 24080 27620 24132
rect 27672 24120 27678 24132
rect 237650 24120 237656 24132
rect 27672 24092 237656 24120
rect 27672 24080 27678 24092
rect 237650 24080 237656 24092
rect 237708 24080 237714 24132
rect 327534 24080 327540 24132
rect 327592 24120 327598 24132
rect 466454 24120 466460 24132
rect 327592 24092 466460 24120
rect 327592 24080 327598 24092
rect 466454 24080 466460 24092
rect 466512 24080 466518 24132
rect 176746 22788 176752 22840
rect 176804 22828 176810 22840
rect 265618 22828 265624 22840
rect 176804 22800 265624 22828
rect 176804 22788 176810 22800
rect 265618 22788 265624 22800
rect 265676 22788 265682 22840
rect 317598 22788 317604 22840
rect 317656 22828 317662 22840
rect 420914 22828 420920 22840
rect 317656 22800 420920 22828
rect 317656 22788 317662 22800
rect 420914 22788 420920 22800
rect 420972 22788 420978 22840
rect 93946 22720 93952 22772
rect 94004 22760 94010 22772
rect 251634 22760 251640 22772
rect 94004 22732 251640 22760
rect 94004 22720 94010 22732
rect 251634 22720 251640 22732
rect 251692 22720 251698 22772
rect 329006 22720 329012 22772
rect 329064 22760 329070 22772
rect 473446 22760 473452 22772
rect 329064 22732 473452 22760
rect 329064 22720 329070 22732
rect 473446 22720 473452 22732
rect 473504 22720 473510 22772
rect 158714 21428 158720 21480
rect 158772 21468 158778 21480
rect 264054 21468 264060 21480
rect 158772 21440 264060 21468
rect 158772 21428 158778 21440
rect 264054 21428 264060 21440
rect 264112 21428 264118 21480
rect 319254 21428 319260 21480
rect 319312 21468 319318 21480
rect 423766 21468 423772 21480
rect 319312 21440 423772 21468
rect 319312 21428 319318 21440
rect 423766 21428 423772 21440
rect 423824 21428 423830 21480
rect 122834 21360 122840 21412
rect 122892 21400 122898 21412
rect 257982 21400 257988 21412
rect 122892 21372 257988 21400
rect 122892 21360 122898 21372
rect 257982 21360 257988 21372
rect 258040 21360 258046 21412
rect 260926 21360 260932 21412
rect 260984 21400 260990 21412
rect 285950 21400 285956 21412
rect 260984 21372 285956 21400
rect 260984 21360 260990 21372
rect 285950 21360 285956 21372
rect 286008 21360 286014 21412
rect 332778 21360 332784 21412
rect 332836 21400 332842 21412
rect 490006 21400 490012 21412
rect 332836 21372 490012 21400
rect 332836 21360 332842 21372
rect 490006 21360 490012 21372
rect 490064 21360 490070 21412
rect 354030 20612 354036 20664
rect 354088 20652 354094 20664
rect 579982 20652 579988 20664
rect 354088 20624 579988 20652
rect 354088 20612 354094 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 297634 20068 297640 20120
rect 297692 20108 297698 20120
rect 318886 20108 318892 20120
rect 297692 20080 318892 20108
rect 297692 20068 297698 20080
rect 318886 20068 318892 20080
rect 318944 20068 318950 20120
rect 144914 20000 144920 20052
rect 144972 20040 144978 20052
rect 261386 20040 261392 20052
rect 144972 20012 261392 20040
rect 144972 20000 144978 20012
rect 261386 20000 261392 20012
rect 261444 20000 261450 20052
rect 306374 20000 306380 20052
rect 306432 20040 306438 20052
rect 365806 20040 365812 20052
rect 306432 20012 365812 20040
rect 306432 20000 306438 20012
rect 365806 20000 365812 20012
rect 365864 20000 365870 20052
rect 30374 19932 30380 19984
rect 30432 19972 30438 19984
rect 238294 19972 238300 19984
rect 30432 19944 238300 19972
rect 30432 19932 30438 19944
rect 238294 19932 238300 19944
rect 238352 19932 238358 19984
rect 258074 19932 258080 19984
rect 258132 19972 258138 19984
rect 285030 19972 285036 19984
rect 258132 19944 285036 19972
rect 258132 19932 258138 19944
rect 285030 19932 285036 19944
rect 285088 19932 285094 19984
rect 318794 19932 318800 19984
rect 318852 19972 318858 19984
rect 425054 19972 425060 19984
rect 318852 19944 425060 19972
rect 318852 19932 318858 19944
rect 425054 19932 425060 19944
rect 425112 19932 425118 19984
rect 118786 18640 118792 18692
rect 118844 18680 118850 18692
rect 255498 18680 255504 18692
rect 118844 18652 255504 18680
rect 118844 18640 118850 18652
rect 255498 18640 255504 18652
rect 255556 18640 255562 18692
rect 320726 18640 320732 18692
rect 320784 18680 320790 18692
rect 432046 18680 432052 18692
rect 320784 18652 432052 18680
rect 320784 18640 320790 18652
rect 432046 18640 432052 18652
rect 432104 18640 432110 18692
rect 49694 18572 49700 18624
rect 49752 18612 49758 18624
rect 242250 18612 242256 18624
rect 49752 18584 242256 18612
rect 49752 18572 49758 18584
rect 242250 18572 242256 18584
rect 242308 18572 242314 18624
rect 242986 18572 242992 18624
rect 243044 18612 243050 18624
rect 281810 18612 281816 18624
rect 243044 18584 281816 18612
rect 243044 18572 243050 18584
rect 281810 18572 281816 18584
rect 281868 18572 281874 18624
rect 296990 18572 296996 18624
rect 297048 18612 297054 18624
rect 316034 18612 316040 18624
rect 297048 18584 316040 18612
rect 297048 18572 297054 18584
rect 316034 18572 316040 18584
rect 316092 18572 316098 18624
rect 332686 18572 332692 18624
rect 332744 18612 332750 18624
rect 492674 18612 492680 18624
rect 332744 18584 492680 18612
rect 332744 18572 332750 18584
rect 492674 18572 492680 18584
rect 492732 18572 492738 18624
rect 226426 17348 226432 17400
rect 226484 17388 226490 17400
rect 278406 17388 278412 17400
rect 226484 17360 278412 17388
rect 226484 17348 226490 17360
rect 278406 17348 278412 17360
rect 278464 17348 278470 17400
rect 85666 17280 85672 17332
rect 85724 17320 85730 17332
rect 248966 17320 248972 17332
rect 85724 17292 248972 17320
rect 85724 17280 85730 17292
rect 248966 17280 248972 17292
rect 249024 17280 249030 17332
rect 311986 17280 311992 17332
rect 312044 17320 312050 17332
rect 393314 17320 393320 17332
rect 312044 17292 393320 17320
rect 312044 17280 312050 17292
rect 393314 17280 393320 17292
rect 393372 17280 393378 17332
rect 2866 17212 2872 17264
rect 2924 17252 2930 17264
rect 231946 17252 231952 17264
rect 2924 17224 231952 17252
rect 2924 17212 2930 17224
rect 231946 17212 231952 17224
rect 232004 17212 232010 17264
rect 301498 17212 301504 17264
rect 301556 17252 301562 17264
rect 339586 17252 339592 17264
rect 301556 17224 339592 17252
rect 301556 17212 301562 17224
rect 339586 17212 339592 17224
rect 339644 17212 339650 17264
rect 355410 17212 355416 17264
rect 355468 17252 355474 17264
rect 576854 17252 576860 17264
rect 355468 17224 576860 17252
rect 355468 17212 355474 17224
rect 576854 17212 576860 17224
rect 576912 17212 576918 17264
rect 205082 15920 205088 15972
rect 205140 15960 205146 15972
rect 274082 15960 274088 15972
rect 205140 15932 274088 15960
rect 205140 15920 205146 15932
rect 274082 15920 274088 15932
rect 274140 15920 274146 15972
rect 339494 15920 339500 15972
rect 339552 15960 339558 15972
rect 523770 15960 523776 15972
rect 339552 15932 523776 15960
rect 339552 15920 339558 15932
rect 523770 15920 523776 15932
rect 523828 15920 523834 15972
rect 69842 15852 69848 15904
rect 69900 15892 69906 15904
rect 246390 15892 246396 15904
rect 69900 15864 246396 15892
rect 69900 15852 69906 15864
rect 246390 15852 246396 15864
rect 246448 15852 246454 15904
rect 299658 15852 299664 15904
rect 299716 15892 299722 15904
rect 328730 15892 328736 15904
rect 299716 15864 328736 15892
rect 299716 15852 299722 15864
rect 328730 15852 328736 15864
rect 328788 15852 328794 15904
rect 346762 15852 346768 15904
rect 346820 15892 346826 15904
rect 560386 15892 560392 15904
rect 346820 15864 560392 15892
rect 346820 15852 346826 15864
rect 560386 15852 560392 15864
rect 560444 15852 560450 15904
rect 298370 14560 298376 14612
rect 298428 14600 298434 14612
rect 324590 14600 324596 14612
rect 298428 14572 324596 14600
rect 298428 14560 298434 14572
rect 324590 14560 324596 14572
rect 324648 14560 324654 14612
rect 116394 14492 116400 14544
rect 116452 14532 116458 14544
rect 255866 14532 255872 14544
rect 116452 14504 255872 14532
rect 116452 14492 116458 14504
rect 255866 14492 255872 14504
rect 255924 14492 255930 14544
rect 277946 14492 277952 14544
rect 278004 14532 278010 14544
rect 289170 14532 289176 14544
rect 278004 14504 289176 14532
rect 278004 14492 278010 14504
rect 289170 14492 289176 14504
rect 289228 14492 289234 14544
rect 317414 14492 317420 14544
rect 317472 14532 317478 14544
rect 415486 14532 415492 14544
rect 317472 14504 415492 14532
rect 317472 14492 317478 14504
rect 415486 14492 415492 14504
rect 415544 14492 415550 14544
rect 53282 14424 53288 14476
rect 53340 14464 53346 14476
rect 242894 14464 242900 14476
rect 53340 14436 242900 14464
rect 53340 14424 53346 14436
rect 242894 14424 242900 14436
rect 242952 14424 242958 14476
rect 251174 14424 251180 14476
rect 251232 14464 251238 14476
rect 283558 14464 283564 14476
rect 251232 14436 283564 14464
rect 251232 14424 251238 14436
rect 283558 14424 283564 14436
rect 283616 14424 283622 14476
rect 305178 14424 305184 14476
rect 305236 14464 305242 14476
rect 357526 14464 357532 14476
rect 305236 14436 357532 14464
rect 305236 14424 305242 14436
rect 357526 14424 357532 14436
rect 357584 14424 357590 14476
rect 364978 14424 364984 14476
rect 365036 14464 365042 14476
rect 568666 14464 568672 14476
rect 365036 14436 568672 14464
rect 365036 14424 365042 14436
rect 568666 14424 568672 14436
rect 568724 14424 568730 14476
rect 270770 13200 270776 13252
rect 270828 13240 270834 13252
rect 287698 13240 287704 13252
rect 270828 13212 287704 13240
rect 270828 13200 270834 13212
rect 287698 13200 287704 13212
rect 287756 13200 287762 13252
rect 309410 13200 309416 13252
rect 309468 13240 309474 13252
rect 376018 13240 376024 13252
rect 309468 13212 376024 13240
rect 309468 13200 309474 13212
rect 376018 13200 376024 13212
rect 376076 13200 376082 13252
rect 190454 13132 190460 13184
rect 190512 13172 190518 13184
rect 271230 13172 271236 13184
rect 190512 13144 271236 13172
rect 190512 13132 190518 13144
rect 271230 13132 271236 13144
rect 271288 13132 271294 13184
rect 320266 13132 320272 13184
rect 320324 13172 320330 13184
rect 429194 13172 429200 13184
rect 320324 13144 429200 13172
rect 320324 13132 320330 13144
rect 429194 13132 429200 13144
rect 429252 13132 429258 13184
rect 91554 13064 91560 13116
rect 91612 13104 91618 13116
rect 250714 13104 250720 13116
rect 91612 13076 250720 13104
rect 91612 13064 91618 13076
rect 250714 13064 250720 13076
rect 250772 13064 250778 13116
rect 252370 13064 252376 13116
rect 252428 13104 252434 13116
rect 283834 13104 283840 13116
rect 252428 13076 283840 13104
rect 252428 13064 252434 13076
rect 283834 13064 283840 13076
rect 283892 13064 283898 13116
rect 302510 13064 302516 13116
rect 302568 13104 302574 13116
rect 345290 13104 345296 13116
rect 302568 13076 345296 13104
rect 302568 13064 302574 13076
rect 345290 13064 345296 13076
rect 345348 13064 345354 13116
rect 363598 13064 363604 13116
rect 363656 13104 363662 13116
rect 551002 13104 551008 13116
rect 363656 13076 551008 13104
rect 363656 13064 363662 13076
rect 551002 13064 551008 13076
rect 551060 13064 551066 13116
rect 75914 11772 75920 11824
rect 75972 11812 75978 11824
rect 247586 11812 247592 11824
rect 75972 11784 247592 11812
rect 75972 11772 75978 11784
rect 247586 11772 247592 11784
rect 247644 11772 247650 11824
rect 264146 11772 264152 11824
rect 264204 11812 264210 11824
rect 286226 11812 286232 11824
rect 264204 11784 286232 11812
rect 264204 11772 264210 11784
rect 286226 11772 286232 11784
rect 286284 11772 286290 11824
rect 309318 11772 309324 11824
rect 309376 11812 309382 11824
rect 379514 11812 379520 11824
rect 309376 11784 379520 11812
rect 309376 11772 309382 11784
rect 379514 11772 379520 11784
rect 379572 11772 379578 11824
rect 71498 11704 71504 11756
rect 71556 11744 71562 11756
rect 246298 11744 246304 11756
rect 71556 11716 246304 11744
rect 71556 11704 71562 11716
rect 246298 11704 246304 11716
rect 246356 11704 246362 11756
rect 247402 11704 247408 11756
rect 247460 11744 247466 11756
rect 283006 11744 283012 11756
rect 247460 11716 283012 11744
rect 247460 11704 247466 11716
rect 283006 11704 283012 11716
rect 283064 11704 283070 11756
rect 301038 11704 301044 11756
rect 301096 11744 301102 11756
rect 338666 11744 338672 11756
rect 301096 11716 338672 11744
rect 301096 11704 301102 11716
rect 338666 11704 338672 11716
rect 338724 11704 338730 11756
rect 352558 11704 352564 11756
rect 352616 11744 352622 11756
rect 533706 11744 533712 11756
rect 352616 11716 533712 11744
rect 352616 11704 352622 11716
rect 533706 11704 533712 11716
rect 533764 11704 533770 11756
rect 160094 11636 160100 11688
rect 160152 11676 160158 11688
rect 161290 11676 161296 11688
rect 160152 11648 161296 11676
rect 160152 11636 160158 11648
rect 161290 11636 161296 11648
rect 161348 11636 161354 11688
rect 176654 11636 176660 11688
rect 176712 11676 176718 11688
rect 177850 11676 177856 11688
rect 176712 11648 177856 11676
rect 176712 11636 176718 11648
rect 177850 11636 177856 11648
rect 177908 11636 177914 11688
rect 184934 11636 184940 11688
rect 184992 11676 184998 11688
rect 186130 11676 186136 11688
rect 184992 11648 186136 11676
rect 184992 11636 184998 11648
rect 186130 11636 186136 11648
rect 186188 11636 186194 11688
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 226334 11636 226340 11688
rect 226392 11676 226398 11688
rect 227530 11676 227536 11688
rect 226392 11648 227536 11676
rect 226392 11636 226398 11648
rect 227530 11636 227536 11648
rect 227588 11636 227594 11688
rect 259454 10412 259460 10464
rect 259512 10452 259518 10464
rect 284478 10452 284484 10464
rect 259512 10424 284484 10452
rect 259512 10412 259518 10424
rect 284478 10412 284484 10424
rect 284536 10412 284542 10464
rect 141234 10344 141240 10396
rect 141292 10384 141298 10396
rect 260098 10384 260104 10396
rect 141292 10356 260104 10384
rect 141292 10344 141298 10356
rect 260098 10344 260104 10356
rect 260156 10344 260162 10396
rect 294690 10344 294696 10396
rect 294748 10384 294754 10396
rect 306374 10384 306380 10396
rect 294748 10356 306380 10384
rect 294748 10344 294754 10356
rect 306374 10344 306380 10356
rect 306432 10344 306438 10396
rect 360838 10344 360844 10396
rect 360896 10384 360902 10396
rect 515490 10384 515496 10396
rect 360896 10356 515496 10384
rect 360896 10344 360902 10356
rect 515490 10344 515496 10356
rect 515548 10344 515554 10396
rect 9674 10276 9680 10328
rect 9732 10316 9738 10328
rect 233970 10316 233976 10328
rect 9732 10288 233976 10316
rect 9732 10276 9738 10288
rect 233970 10276 233976 10288
rect 234028 10276 234034 10328
rect 234614 10276 234620 10328
rect 234672 10316 234678 10328
rect 279510 10316 279516 10328
rect 234672 10288 279516 10316
rect 234672 10276 234678 10288
rect 279510 10276 279516 10288
rect 279568 10276 279574 10328
rect 305730 10276 305736 10328
rect 305788 10316 305794 10328
rect 321646 10316 321652 10328
rect 305788 10288 321652 10316
rect 305788 10276 305794 10288
rect 321646 10276 321652 10288
rect 321704 10276 321710 10328
rect 341150 10276 341156 10328
rect 341208 10316 341214 10328
rect 532050 10316 532056 10328
rect 341208 10288 532056 10316
rect 341208 10276 341214 10288
rect 532050 10276 532056 10288
rect 532108 10276 532114 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 254670 9052 254676 9104
rect 254728 9092 254734 9104
rect 280798 9092 280804 9104
rect 254728 9064 280804 9092
rect 254728 9052 254734 9064
rect 280798 9052 280804 9064
rect 280856 9052 280862 9104
rect 293770 9052 293776 9104
rect 293828 9092 293834 9104
rect 300762 9092 300768 9104
rect 293828 9064 300768 9092
rect 293828 9052 293834 9064
rect 300762 9052 300768 9064
rect 300820 9052 300826 9104
rect 137646 8984 137652 9036
rect 137704 9024 137710 9036
rect 224218 9024 224224 9036
rect 137704 8996 224224 9024
rect 137704 8984 137710 8996
rect 224218 8984 224224 8996
rect 224276 8984 224282 9036
rect 238110 8984 238116 9036
rect 238168 9024 238174 9036
rect 280614 9024 280620 9036
rect 238168 8996 280620 9024
rect 238168 8984 238174 8996
rect 280614 8984 280620 8996
rect 280672 8984 280678 9036
rect 298094 8984 298100 9036
rect 298152 9024 298158 9036
rect 326798 9024 326804 9036
rect 298152 8996 326804 9024
rect 298152 8984 298158 8996
rect 326798 8984 326804 8996
rect 326856 8984 326862 9036
rect 355318 8984 355324 9036
rect 355376 9024 355382 9036
rect 505370 9024 505376 9036
rect 355376 8996 505376 9024
rect 355376 8984 355382 8996
rect 505370 8984 505376 8996
rect 505428 8984 505434 9036
rect 38378 8916 38384 8968
rect 38436 8956 38442 8968
rect 239674 8956 239680 8968
rect 38436 8928 239680 8956
rect 38436 8916 38442 8928
rect 239674 8916 239680 8928
rect 239732 8916 239738 8968
rect 246390 8916 246396 8968
rect 246448 8956 246454 8968
rect 282546 8956 282552 8968
rect 246448 8928 282552 8956
rect 246448 8916 246454 8928
rect 282546 8916 282552 8928
rect 282604 8916 282610 8968
rect 299474 8916 299480 8968
rect 299532 8956 299538 8968
rect 327994 8956 328000 8968
rect 299532 8928 328000 8956
rect 299532 8916 299538 8928
rect 327994 8916 328000 8928
rect 328052 8916 328058 8968
rect 336826 8916 336832 8968
rect 336884 8956 336890 8968
rect 514754 8956 514760 8968
rect 336884 8928 514760 8956
rect 336884 8916 336890 8928
rect 514754 8916 514760 8928
rect 514812 8916 514818 8968
rect 307110 8236 307116 8288
rect 307168 8276 307174 8288
rect 309042 8276 309048 8288
rect 307168 8248 309048 8276
rect 307168 8236 307174 8248
rect 309042 8236 309048 8248
rect 309100 8236 309106 8288
rect 241698 7760 241704 7812
rect 241756 7800 241762 7812
rect 273898 7800 273904 7812
rect 241756 7772 273904 7800
rect 241756 7760 241762 7772
rect 273898 7760 273904 7772
rect 273956 7760 273962 7812
rect 218146 7692 218152 7744
rect 218204 7732 218210 7744
rect 225598 7732 225604 7744
rect 218204 7704 225604 7732
rect 218204 7692 218210 7704
rect 225598 7692 225604 7704
rect 225656 7692 225662 7744
rect 242894 7692 242900 7744
rect 242952 7732 242958 7744
rect 281902 7732 281908 7744
rect 242952 7704 281908 7732
rect 242952 7692 242958 7704
rect 281902 7692 281908 7704
rect 281960 7692 281966 7744
rect 92750 7624 92756 7676
rect 92808 7664 92814 7676
rect 250438 7664 250444 7676
rect 92808 7636 250444 7664
rect 92808 7624 92814 7636
rect 250438 7624 250444 7636
rect 250496 7624 250502 7676
rect 296162 7624 296168 7676
rect 296220 7664 296226 7676
rect 312630 7664 312636 7676
rect 296220 7636 312636 7664
rect 296220 7624 296226 7636
rect 312630 7624 312636 7636
rect 312688 7624 312694 7676
rect 359458 7624 359464 7676
rect 359516 7664 359522 7676
rect 501782 7664 501788 7676
rect 359516 7636 501788 7664
rect 359516 7624 359522 7636
rect 501782 7624 501788 7636
rect 501840 7624 501846 7676
rect 51350 7556 51356 7608
rect 51408 7596 51414 7608
rect 221458 7596 221464 7608
rect 51408 7568 221464 7596
rect 51408 7556 51414 7568
rect 221458 7556 221464 7568
rect 221516 7556 221522 7608
rect 233418 7556 233424 7608
rect 233476 7596 233482 7608
rect 279142 7596 279148 7608
rect 233476 7568 279148 7596
rect 233476 7556 233482 7568
rect 279142 7556 279148 7568
rect 279200 7556 279206 7608
rect 297358 7556 297364 7608
rect 297416 7596 297422 7608
rect 320910 7596 320916 7608
rect 297416 7568 320916 7596
rect 297416 7556 297422 7568
rect 320910 7556 320916 7568
rect 320968 7556 320974 7608
rect 335354 7556 335360 7608
rect 335412 7596 335418 7608
rect 507670 7596 507676 7608
rect 335412 7568 507676 7596
rect 335412 7556 335418 7568
rect 507670 7556 507676 7568
rect 507728 7556 507734 7608
rect 281902 6876 281908 6928
rect 281960 6916 281966 6928
rect 289078 6916 289084 6928
rect 281960 6888 289084 6916
rect 281960 6876 281966 6888
rect 289078 6876 289084 6888
rect 289136 6876 289142 6928
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 229738 6848 229744 6860
rect 3476 6820 229744 6848
rect 3476 6808 3482 6820
rect 229738 6808 229744 6820
rect 229796 6808 229802 6860
rect 353938 6808 353944 6860
rect 353996 6848 354002 6860
rect 580166 6848 580172 6860
rect 353996 6820 580172 6848
rect 353996 6808 354002 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 239306 6332 239312 6384
rect 239364 6372 239370 6384
rect 268378 6372 268384 6384
rect 239364 6344 268384 6372
rect 239364 6332 239370 6344
rect 268378 6332 268384 6344
rect 268436 6332 268442 6384
rect 276014 6332 276020 6384
rect 276072 6372 276078 6384
rect 284938 6372 284944 6384
rect 276072 6344 284944 6372
rect 276072 6332 276078 6344
rect 284938 6332 284944 6344
rect 284996 6332 285002 6384
rect 253474 6264 253480 6316
rect 253532 6304 253538 6316
rect 283282 6304 283288 6316
rect 253532 6276 283288 6304
rect 253532 6264 253538 6276
rect 283282 6264 283288 6276
rect 283340 6264 283346 6316
rect 296898 6264 296904 6316
rect 296956 6304 296962 6316
rect 318518 6304 318524 6316
rect 296956 6276 318524 6304
rect 296956 6264 296962 6276
rect 318518 6264 318524 6276
rect 318576 6264 318582 6316
rect 240502 6196 240508 6248
rect 240560 6236 240566 6248
rect 278130 6236 278136 6248
rect 240560 6208 278136 6236
rect 240560 6196 240566 6208
rect 278130 6196 278136 6208
rect 278188 6196 278194 6248
rect 303706 6196 303712 6248
rect 303764 6236 303770 6248
rect 351638 6236 351644 6248
rect 303764 6208 351644 6236
rect 303764 6196 303770 6208
rect 351638 6196 351644 6208
rect 351696 6196 351702 6248
rect 78582 6128 78588 6180
rect 78640 6168 78646 6180
rect 247494 6168 247500 6180
rect 78640 6140 247500 6168
rect 78640 6128 78646 6140
rect 247494 6128 247500 6140
rect 247552 6128 247558 6180
rect 248782 6128 248788 6180
rect 248840 6168 248846 6180
rect 282178 6168 282184 6180
rect 248840 6140 282184 6168
rect 248840 6128 248846 6140
rect 282178 6128 282184 6140
rect 282236 6128 282242 6180
rect 313458 6128 313464 6180
rect 313516 6168 313522 6180
rect 397730 6168 397736 6180
rect 313516 6140 397736 6168
rect 313516 6128 313522 6140
rect 397730 6128 397736 6140
rect 397788 6128 397794 6180
rect 295886 6060 295892 6112
rect 295944 6100 295950 6112
rect 313826 6100 313832 6112
rect 295944 6072 313832 6100
rect 295944 6060 295950 6072
rect 313826 6060 313832 6072
rect 313884 6060 313890 6112
rect 293494 5448 293500 5500
rect 293552 5488 293558 5500
rect 299658 5488 299664 5500
rect 293552 5460 299664 5488
rect 293552 5448 293558 5460
rect 299658 5448 299664 5460
rect 299716 5448 299722 5500
rect 249978 4972 249984 5024
rect 250036 5012 250042 5024
rect 275278 5012 275284 5024
rect 250036 4984 275284 5012
rect 250036 4972 250042 4984
rect 275278 4972 275284 4984
rect 275336 4972 275342 5024
rect 237006 4904 237012 4956
rect 237064 4944 237070 4956
rect 269758 4944 269764 4956
rect 237064 4916 269764 4944
rect 237064 4904 237070 4916
rect 269758 4904 269764 4916
rect 269816 4904 269822 4956
rect 272426 4904 272432 4956
rect 272484 4944 272490 4956
rect 287974 4944 287980 4956
rect 272484 4916 287980 4944
rect 272484 4904 272490 4916
rect 287974 4904 287980 4916
rect 288032 4904 288038 4956
rect 295702 4904 295708 4956
rect 295760 4944 295766 4956
rect 310238 4944 310244 4956
rect 295760 4916 310244 4944
rect 295760 4904 295766 4916
rect 310238 4904 310244 4916
rect 310296 4904 310302 4956
rect 168466 4836 168472 4888
rect 168524 4876 168530 4888
rect 228358 4876 228364 4888
rect 168524 4848 228364 4876
rect 168524 4836 168530 4848
rect 228358 4836 228364 4848
rect 228416 4836 228422 4888
rect 235810 4836 235816 4888
rect 235868 4876 235874 4888
rect 278038 4876 278044 4888
rect 235868 4848 278044 4876
rect 235868 4836 235874 4848
rect 278038 4836 278044 4848
rect 278096 4836 278102 4888
rect 295426 4836 295432 4888
rect 295484 4876 295490 4888
rect 311434 4876 311440 4888
rect 295484 4848 311440 4876
rect 295484 4836 295490 4848
rect 311434 4836 311440 4848
rect 311492 4836 311498 4888
rect 334158 4836 334164 4888
rect 334216 4876 334222 4888
rect 334216 4848 335354 4876
rect 334216 4836 334222 4848
rect 34790 4768 34796 4820
rect 34848 4808 34854 4820
rect 239214 4808 239220 4820
rect 34848 4780 239220 4808
rect 34848 4768 34854 4780
rect 239214 4768 239220 4780
rect 239272 4768 239278 4820
rect 245194 4768 245200 4820
rect 245252 4808 245258 4820
rect 282270 4808 282276 4820
rect 245252 4780 282276 4808
rect 245252 4768 245258 4780
rect 282270 4768 282276 4780
rect 282328 4768 282334 4820
rect 299566 4768 299572 4820
rect 299624 4808 299630 4820
rect 330386 4808 330392 4820
rect 299624 4780 330392 4808
rect 299624 4768 299630 4780
rect 330386 4768 330392 4780
rect 330444 4768 330450 4820
rect 335326 4808 335354 4848
rect 356698 4836 356704 4888
rect 356756 4876 356762 4888
rect 484026 4876 484032 4888
rect 356756 4848 484032 4876
rect 356756 4836 356762 4848
rect 484026 4836 484032 4848
rect 484084 4836 484090 4888
rect 497090 4808 497096 4820
rect 335326 4780 497096 4808
rect 497090 4768 497096 4780
rect 497148 4768 497154 4820
rect 311158 4428 311164 4480
rect 311216 4468 311222 4480
rect 317322 4468 317328 4480
rect 311216 4440 317328 4468
rect 311216 4428 311222 4440
rect 317322 4428 317328 4440
rect 317380 4428 317386 4480
rect 274818 4292 274824 4344
rect 274876 4332 274882 4344
rect 279418 4332 279424 4344
rect 274876 4304 279424 4332
rect 274876 4292 274882 4304
rect 279418 4292 279424 4304
rect 279476 4292 279482 4344
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 193214 4156 193220 4208
rect 193272 4196 193278 4208
rect 194410 4196 194416 4208
rect 193272 4168 194416 4196
rect 193272 4156 193278 4168
rect 194410 4156 194416 4168
rect 194468 4156 194474 4208
rect 218054 4156 218060 4208
rect 218112 4196 218118 4208
rect 219250 4196 219256 4208
rect 218112 4168 219256 4196
rect 218112 4156 218118 4168
rect 219250 4156 219256 4168
rect 219308 4156 219314 4208
rect 307018 4156 307024 4208
rect 307076 4196 307082 4208
rect 307938 4196 307944 4208
rect 307076 4168 307944 4196
rect 307076 4156 307082 4168
rect 307938 4156 307944 4168
rect 307996 4156 308002 4208
rect 319438 4156 319444 4208
rect 319496 4196 319502 4208
rect 324314 4196 324320 4208
rect 319496 4168 324320 4196
rect 319496 4156 319502 4168
rect 324314 4156 324320 4168
rect 324372 4156 324378 4208
rect 331858 4156 331864 4208
rect 331916 4196 331922 4208
rect 335078 4196 335084 4208
rect 331916 4168 335084 4196
rect 331916 4156 331922 4168
rect 335078 4156 335084 4168
rect 335136 4156 335142 4208
rect 485038 4156 485044 4208
rect 485096 4196 485102 4208
rect 487614 4196 487620 4208
rect 485096 4168 487620 4196
rect 485096 4156 485102 4168
rect 487614 4156 487620 4168
rect 487672 4156 487678 4208
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 240686 4128 240692 4140
rect 43128 4100 240692 4128
rect 43128 4088 43134 4100
rect 240686 4088 240692 4100
rect 240744 4088 240750 4140
rect 284294 4088 284300 4140
rect 284352 4128 284358 4140
rect 290366 4128 290372 4140
rect 284352 4100 290372 4128
rect 284352 4088 284358 4100
rect 290366 4088 290372 4100
rect 290424 4088 290430 4140
rect 292666 4088 292672 4140
rect 292724 4128 292730 4140
rect 294874 4128 294880 4140
rect 292724 4100 294880 4128
rect 292724 4088 292730 4100
rect 294874 4088 294880 4100
rect 294932 4088 294938 4140
rect 324682 4088 324688 4140
rect 324740 4128 324746 4140
rect 450906 4128 450912 4140
rect 324740 4100 450912 4128
rect 324740 4088 324746 4100
rect 450906 4088 450912 4100
rect 450964 4088 450970 4140
rect 39574 4020 39580 4072
rect 39632 4060 39638 4072
rect 241422 4060 241428 4072
rect 39632 4032 241428 4060
rect 39632 4020 39638 4032
rect 241422 4020 241428 4032
rect 241480 4020 241486 4072
rect 283098 4020 283104 4072
rect 283156 4060 283162 4072
rect 290182 4060 290188 4072
rect 283156 4032 290188 4060
rect 283156 4020 283162 4032
rect 290182 4020 290188 4032
rect 290240 4020 290246 4072
rect 292850 4020 292856 4072
rect 292908 4060 292914 4072
rect 296070 4060 296076 4072
rect 292908 4032 296076 4060
rect 292908 4020 292914 4032
rect 296070 4020 296076 4032
rect 296128 4020 296134 4072
rect 324406 4020 324412 4072
rect 324464 4060 324470 4072
rect 454494 4060 454500 4072
rect 324464 4032 454500 4060
rect 324464 4020 324470 4032
rect 454494 4020 454500 4032
rect 454552 4020 454558 4072
rect 35986 3952 35992 4004
rect 36044 3992 36050 4004
rect 238754 3992 238760 4004
rect 36044 3964 238760 3992
rect 36044 3952 36050 3964
rect 238754 3952 238760 3964
rect 238812 3952 238818 4004
rect 292758 3952 292764 4004
rect 292816 3992 292822 4004
rect 297266 3992 297272 4004
rect 292816 3964 297272 3992
rect 292816 3952 292822 3964
rect 297266 3952 297272 3964
rect 297324 3952 297330 4004
rect 326062 3952 326068 4004
rect 326120 3992 326126 4004
rect 458082 3992 458088 4004
rect 326120 3964 458088 3992
rect 326120 3952 326126 3964
rect 458082 3952 458088 3964
rect 458140 3952 458146 4004
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 238018 3924 238024 3936
rect 32456 3896 238024 3924
rect 32456 3884 32462 3896
rect 238018 3884 238024 3896
rect 238076 3884 238082 3936
rect 279510 3884 279516 3936
rect 279568 3924 279574 3936
rect 289354 3924 289360 3936
rect 279568 3896 289360 3924
rect 279568 3884 279574 3896
rect 289354 3884 289360 3896
rect 289412 3884 289418 3936
rect 293218 3884 293224 3936
rect 293276 3924 293282 3936
rect 298462 3924 298468 3936
rect 293276 3896 298468 3924
rect 293276 3884 293282 3896
rect 298462 3884 298468 3896
rect 298520 3884 298526 3936
rect 326338 3884 326344 3936
rect 326396 3924 326402 3936
rect 461578 3924 461584 3936
rect 326396 3896 461584 3924
rect 326396 3884 326402 3896
rect 461578 3884 461584 3896
rect 461636 3884 461642 3936
rect 28902 3816 28908 3868
rect 28960 3856 28966 3868
rect 237834 3856 237840 3868
rect 28960 3828 237840 3856
rect 28960 3816 28966 3828
rect 237834 3816 237840 3828
rect 237892 3816 237898 3868
rect 277118 3816 277124 3868
rect 277176 3856 277182 3868
rect 288618 3856 288624 3868
rect 277176 3828 288624 3856
rect 277176 3816 277182 3828
rect 288618 3816 288624 3828
rect 288676 3816 288682 3868
rect 293954 3816 293960 3868
rect 294012 3856 294018 3868
rect 301958 3856 301964 3868
rect 294012 3828 301964 3856
rect 294012 3816 294018 3828
rect 301958 3816 301964 3828
rect 302016 3816 302022 3868
rect 327074 3816 327080 3868
rect 327132 3856 327138 3868
rect 465166 3856 465172 3868
rect 327132 3828 465172 3856
rect 327132 3816 327138 3828
rect 465166 3816 465172 3828
rect 465224 3816 465230 3868
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 236914 3788 236920 3800
rect 25372 3760 236920 3788
rect 25372 3748 25378 3760
rect 236914 3748 236920 3760
rect 236972 3748 236978 3800
rect 273622 3748 273628 3800
rect 273680 3788 273686 3800
rect 287882 3788 287888 3800
rect 273680 3760 287888 3788
rect 273680 3748 273686 3760
rect 287882 3748 287888 3760
rect 287940 3748 287946 3800
rect 328454 3748 328460 3800
rect 328512 3788 328518 3800
rect 468662 3788 468668 3800
rect 328512 3760 468668 3788
rect 328512 3748 328518 3760
rect 468662 3748 468668 3760
rect 468720 3748 468726 3800
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 236822 3720 236828 3732
rect 24268 3692 236828 3720
rect 24268 3680 24274 3692
rect 236822 3680 236828 3692
rect 236880 3680 236886 3732
rect 267734 3680 267740 3732
rect 267792 3720 267798 3732
rect 268470 3720 268476 3732
rect 267792 3692 268476 3720
rect 267792 3680 267798 3692
rect 268470 3680 268476 3692
rect 268528 3680 268534 3732
rect 270034 3680 270040 3732
rect 270092 3720 270098 3732
rect 287146 3720 287152 3732
rect 270092 3692 287152 3720
rect 270092 3680 270098 3692
rect 287146 3680 287152 3692
rect 287204 3680 287210 3732
rect 328546 3680 328552 3732
rect 328604 3720 328610 3732
rect 472250 3720 472256 3732
rect 328604 3692 472256 3720
rect 328604 3680 328610 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 10318 3652 10324 3664
rect 6886 3624 10324 3652
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 4798 3516 4804 3528
rect 624 3488 4804 3516
rect 624 3476 630 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6886 3516 6914 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 235994 3652 236000 3664
rect 19484 3624 236000 3652
rect 19484 3612 19490 3624
rect 235994 3612 236000 3624
rect 236052 3612 236058 3664
rect 266538 3612 266544 3664
rect 266596 3652 266602 3664
rect 286410 3652 286416 3664
rect 266596 3624 286416 3652
rect 266596 3612 266602 3624
rect 286410 3612 286416 3624
rect 286468 3612 286474 3664
rect 329834 3612 329840 3664
rect 329892 3652 329898 3664
rect 475746 3652 475752 3664
rect 329892 3624 475752 3652
rect 329892 3612 329898 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 7558 3544 7564 3596
rect 7616 3544 7622 3596
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 236270 3584 236276 3596
rect 20680 3556 236276 3584
rect 20680 3544 20686 3556
rect 236270 3544 236276 3556
rect 236328 3544 236334 3596
rect 262950 3544 262956 3596
rect 263008 3584 263014 3596
rect 285674 3584 285680 3596
rect 263008 3556 285680 3584
rect 263008 3544 263014 3556
rect 285674 3544 285680 3556
rect 285732 3544 285738 3596
rect 286594 3544 286600 3596
rect 286652 3584 286658 3596
rect 290090 3584 290096 3596
rect 286652 3556 290096 3584
rect 286652 3544 286658 3556
rect 290090 3544 290096 3556
rect 290148 3544 290154 3596
rect 291562 3544 291568 3596
rect 291620 3584 291626 3596
rect 293678 3584 293684 3596
rect 291620 3556 293684 3584
rect 291620 3544 291626 3556
rect 293678 3544 293684 3556
rect 293736 3544 293742 3596
rect 321738 3544 321744 3596
rect 321796 3584 321802 3596
rect 321796 3556 321876 3584
rect 321796 3544 321802 3556
rect 5316 3488 6914 3516
rect 5316 3476 5322 3488
rect 1670 3272 1676 3324
rect 1728 3312 1734 3324
rect 7576 3312 7604 3544
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 235074 3516 235080 3528
rect 15988 3488 235080 3516
rect 15988 3476 15994 3488
rect 235074 3476 235080 3488
rect 235132 3476 235138 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260650 3516 260656 3528
rect 259512 3488 260656 3516
rect 259512 3476 259518 3488
rect 260650 3476 260656 3488
rect 260708 3476 260714 3528
rect 285398 3476 285404 3528
rect 285456 3516 285462 3528
rect 290550 3516 290556 3528
rect 285456 3488 290556 3516
rect 285456 3476 285462 3488
rect 290550 3476 290556 3488
rect 290608 3476 290614 3528
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 233602 3448 233608 3460
rect 11204 3420 233608 3448
rect 11204 3408 11210 3420
rect 233602 3408 233608 3420
rect 233660 3408 233666 3460
rect 255866 3408 255872 3460
rect 255924 3448 255930 3460
rect 285214 3448 285220 3460
rect 255924 3420 285220 3448
rect 255924 3408 255930 3420
rect 285214 3408 285220 3420
rect 285272 3408 285278 3460
rect 292022 3408 292028 3460
rect 292080 3448 292086 3460
rect 292574 3448 292580 3460
rect 292080 3420 292580 3448
rect 292080 3408 292086 3420
rect 292574 3408 292580 3420
rect 292632 3408 292638 3460
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 241514 3380 241520 3392
rect 46716 3352 241520 3380
rect 46716 3340 46722 3352
rect 241514 3340 241520 3352
rect 241572 3340 241578 3392
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 285306 3380 285312 3392
rect 259512 3352 285312 3380
rect 259512 3340 259518 3352
rect 285306 3340 285312 3352
rect 285364 3340 285370 3392
rect 294230 3340 294236 3392
rect 294288 3380 294294 3392
rect 305546 3380 305552 3392
rect 294288 3352 305552 3380
rect 294288 3340 294294 3352
rect 305546 3340 305552 3352
rect 305604 3340 305610 3392
rect 1728 3284 7604 3312
rect 1728 3272 1734 3284
rect 60734 3272 60740 3324
rect 60792 3312 60798 3324
rect 61654 3312 61660 3324
rect 60792 3284 61660 3312
rect 60792 3272 60798 3284
rect 61654 3272 61660 3284
rect 61712 3272 61718 3324
rect 85574 3272 85580 3324
rect 85632 3312 85638 3324
rect 86494 3312 86500 3324
rect 85632 3284 86500 3312
rect 85632 3272 85638 3284
rect 86494 3272 86500 3284
rect 86552 3272 86558 3324
rect 110414 3272 110420 3324
rect 110472 3312 110478 3324
rect 111610 3312 111616 3324
rect 110472 3284 111616 3312
rect 110472 3272 110478 3284
rect 111610 3272 111616 3284
rect 111668 3272 111674 3324
rect 118694 3272 118700 3324
rect 118752 3312 118758 3324
rect 119890 3312 119896 3324
rect 118752 3284 119896 3312
rect 118752 3272 118758 3284
rect 119890 3272 119896 3284
rect 119948 3272 119954 3324
rect 255774 3312 255780 3324
rect 120092 3284 255780 3312
rect 117590 3204 117596 3256
rect 117648 3244 117654 3256
rect 120092 3244 120120 3284
rect 255774 3272 255780 3284
rect 255832 3272 255838 3324
rect 280706 3272 280712 3324
rect 280764 3312 280770 3324
rect 289630 3312 289636 3324
rect 280764 3284 289636 3312
rect 280764 3272 280770 3284
rect 289630 3272 289636 3284
rect 289688 3272 289694 3324
rect 290182 3272 290188 3324
rect 290240 3312 290246 3324
rect 291654 3312 291660 3324
rect 290240 3284 291660 3312
rect 290240 3272 290246 3284
rect 291654 3272 291660 3284
rect 291712 3272 291718 3324
rect 117648 3216 120120 3244
rect 117648 3204 117654 3216
rect 121086 3204 121092 3256
rect 121144 3244 121150 3256
rect 257246 3244 257252 3256
rect 121144 3216 257252 3244
rect 121144 3204 121150 3216
rect 257246 3204 257252 3216
rect 257304 3204 257310 3256
rect 321848 3244 321876 3556
rect 351178 3544 351184 3596
rect 351236 3584 351242 3596
rect 582190 3584 582196 3596
rect 351236 3556 582196 3584
rect 351236 3544 351242 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 330202 3476 330208 3528
rect 330260 3516 330266 3528
rect 479334 3516 479340 3528
rect 330260 3488 479340 3516
rect 330260 3476 330266 3488
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 563698 3476 563704 3528
rect 563756 3516 563762 3528
rect 564434 3516 564440 3528
rect 563756 3488 564440 3516
rect 563756 3476 563762 3488
rect 564434 3476 564440 3488
rect 564492 3476 564498 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 572714 3516 572720 3528
rect 572036 3488 572720 3516
rect 572036 3476 572042 3488
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 349246 3408 349252 3460
rect 349304 3448 349310 3460
rect 350442 3448 350448 3460
rect 349304 3420 350448 3448
rect 349304 3408 349310 3420
rect 350442 3408 350448 3420
rect 350500 3408 350506 3460
rect 350902 3408 350908 3460
rect 350960 3448 350966 3460
rect 580994 3448 581000 3460
rect 350960 3420 581000 3448
rect 350960 3408 350966 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 323394 3340 323400 3392
rect 323452 3380 323458 3392
rect 447410 3380 447416 3392
rect 323452 3352 447416 3380
rect 323452 3340 323458 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 322934 3272 322940 3324
rect 322992 3312 322998 3324
rect 443822 3312 443828 3324
rect 322992 3284 443828 3312
rect 322992 3272 322998 3284
rect 443822 3272 443828 3284
rect 443880 3272 443886 3324
rect 440234 3244 440240 3256
rect 321848 3216 440240 3244
rect 440234 3204 440240 3216
rect 440292 3204 440298 3256
rect 440326 3204 440332 3256
rect 440384 3244 440390 3256
rect 441522 3244 441528 3256
rect 440384 3216 441528 3244
rect 440384 3204 440390 3216
rect 441522 3204 441528 3216
rect 441580 3204 441586 3256
rect 168374 3136 168380 3188
rect 168432 3176 168438 3188
rect 169570 3176 169576 3188
rect 168432 3148 169576 3176
rect 168432 3136 168438 3148
rect 169570 3136 169576 3148
rect 169628 3136 169634 3188
rect 288986 3136 288992 3188
rect 289044 3176 289050 3188
rect 291286 3176 291292 3188
rect 289044 3148 291292 3176
rect 289044 3136 289050 3148
rect 291286 3136 291292 3148
rect 291344 3136 291350 3188
rect 357526 3136 357532 3188
rect 357584 3176 357590 3188
rect 358722 3176 358728 3188
rect 357584 3148 358728 3176
rect 357584 3136 357590 3148
rect 358722 3136 358728 3148
rect 358780 3136 358786 3188
rect 374086 3136 374092 3188
rect 374144 3176 374150 3188
rect 375282 3176 375288 3188
rect 374144 3148 375288 3176
rect 374144 3136 374150 3148
rect 375282 3136 375288 3148
rect 375340 3136 375346 3188
rect 382366 3136 382372 3188
rect 382424 3176 382430 3188
rect 383562 3176 383568 3188
rect 382424 3148 383568 3176
rect 382424 3136 382430 3148
rect 383562 3136 383568 3148
rect 383620 3136 383626 3188
rect 398926 3136 398932 3188
rect 398984 3176 398990 3188
rect 400122 3176 400128 3188
rect 398984 3148 400128 3176
rect 398984 3136 398990 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 407114 3136 407120 3188
rect 407172 3176 407178 3188
rect 408402 3176 408408 3188
rect 407172 3148 408408 3176
rect 407172 3136 407178 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 415394 3136 415400 3188
rect 415452 3176 415458 3188
rect 416682 3176 416688 3188
rect 415452 3148 416688 3176
rect 415452 3136 415458 3148
rect 416682 3136 416688 3148
rect 416740 3136 416746 3188
rect 423766 3136 423772 3188
rect 423824 3176 423830 3188
rect 424962 3176 424968 3188
rect 423824 3148 424968 3176
rect 423824 3136 423830 3148
rect 424962 3136 424968 3148
rect 425020 3136 425026 3188
rect 431954 3136 431960 3188
rect 432012 3176 432018 3188
rect 433242 3176 433248 3188
rect 432012 3148 433248 3176
rect 432012 3136 432018 3148
rect 433242 3136 433248 3148
rect 433300 3136 433306 3188
rect 287790 3068 287796 3120
rect 287848 3108 287854 3120
rect 291194 3108 291200 3120
rect 287848 3080 291200 3108
rect 287848 3068 287854 3080
rect 291194 3068 291200 3080
rect 291252 3068 291258 3120
rect 340874 2728 340880 2780
rect 340932 2768 340938 2780
rect 342162 2768 342168 2780
rect 340932 2740 342168 2768
rect 340932 2728 340938 2740
rect 342162 2728 342168 2740
rect 342220 2728 342226 2780
rect 365714 1504 365720 1556
rect 365772 1544 365778 1556
rect 367002 1544 367008 1556
rect 365772 1516 367008 1544
rect 365772 1504 365778 1516
rect 367002 1504 367008 1516
rect 367060 1504 367066 1556
rect 390554 1504 390560 1556
rect 390612 1544 390618 1556
rect 391842 1544 391848 1556
rect 390612 1516 391848 1544
rect 390612 1504 390618 1516
rect 391842 1504 391848 1516
rect 391900 1504 391906 1556
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 309140 700884 309192 700936
rect 364984 700884 365036 700936
rect 313280 700816 313332 700868
rect 397460 700816 397512 700868
rect 317420 700748 317472 700800
rect 413652 700748 413704 700800
rect 322940 700680 322992 700732
rect 429844 700680 429896 700732
rect 327080 700612 327132 700664
rect 462320 700612 462372 700664
rect 331312 700544 331364 700596
rect 478512 700544 478564 700596
rect 335360 700476 335412 700528
rect 494796 700476 494848 700528
rect 340880 700408 340932 700460
rect 527180 700408 527232 700460
rect 300860 700340 300912 700392
rect 332508 700340 332560 700392
rect 345020 700340 345072 700392
rect 543464 700340 543516 700392
rect 267648 700272 267700 700324
rect 279424 700272 279476 700324
rect 295340 700272 295392 700324
rect 300124 700272 300176 700324
rect 305000 700272 305052 700324
rect 348792 700272 348844 700324
rect 349160 700272 349212 700324
rect 559656 700272 559708 700324
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 353944 683136 353996 683188
rect 579620 683136 579672 683188
rect 360844 670692 360896 670744
rect 580172 670692 580224 670744
rect 367744 643084 367796 643136
rect 580172 643084 580224 643136
rect 3332 632068 3384 632120
rect 32404 632068 32456 632120
rect 374644 630640 374696 630692
rect 579988 630640 580040 630692
rect 3332 618264 3384 618316
rect 22744 618264 22796 618316
rect 381544 616836 381596 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 14464 605820 14516 605872
rect 3148 579776 3200 579828
rect 7564 579776 7616 579828
rect 359464 563048 359516 563100
rect 580172 563048 580224 563100
rect 364984 536800 365036 536852
rect 580172 536800 580224 536852
rect 2964 527144 3016 527196
rect 43444 527144 43496 527196
rect 373264 524424 373316 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 25504 514768 25556 514820
rect 356704 510620 356756 510672
rect 580172 510620 580224 510672
rect 3240 500964 3292 501016
rect 17224 500964 17276 501016
rect 3332 475192 3384 475244
rect 8944 475192 8996 475244
rect 355324 456764 355376 456816
rect 580172 456764 580224 456816
rect 371884 430584 371936 430636
rect 580172 430584 580224 430636
rect 2964 422288 3016 422340
rect 31024 422288 31076 422340
rect 378784 418140 378836 418192
rect 580172 418140 580224 418192
rect 3332 409844 3384 409896
rect 26884 409844 26936 409896
rect 363604 404336 363656 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 18604 397468 18656 397520
rect 3332 371220 3384 371272
rect 10324 371220 10376 371272
rect 354036 364352 354088 364404
rect 580172 364352 580224 364404
rect 369124 324300 369176 324352
rect 579988 324300 580040 324352
rect 3148 318792 3200 318844
rect 221464 318792 221516 318844
rect 377404 311856 377456 311908
rect 579804 311856 579856 311908
rect 3332 304988 3384 305040
rect 28264 304988 28316 305040
rect 442264 298120 442316 298172
rect 580172 298120 580224 298172
rect 3332 292544 3384 292596
rect 21364 292544 21416 292596
rect 3240 266364 3292 266416
rect 13084 266364 13136 266416
rect 218060 263508 218112 263560
rect 278596 263508 278648 263560
rect 201500 263440 201552 263492
rect 274180 263440 274232 263492
rect 169760 263372 169812 263424
rect 269764 263372 269816 263424
rect 153200 263304 153252 263356
rect 265348 263304 265400 263356
rect 136640 263236 136692 263288
rect 260840 263236 260892 263288
rect 104900 263168 104952 263220
rect 256424 263168 256476 263220
rect 88340 263100 88392 263152
rect 252008 263100 252060 263152
rect 71780 263032 71832 263084
rect 247500 263032 247552 263084
rect 40040 262964 40092 263016
rect 243084 262964 243136 263016
rect 282920 262964 282972 263016
rect 291936 262964 291988 263016
rect 23480 262896 23532 262948
rect 238668 262896 238720 262948
rect 279424 262896 279476 262948
rect 287520 262896 287572 262948
rect 6920 262828 6972 262880
rect 234252 262828 234304 262880
rect 234620 262828 234672 262880
rect 283104 262828 283156 262880
rect 4804 259360 4856 259412
rect 229100 259360 229152 259412
rect 354312 259360 354364 259412
rect 580264 259360 580316 259412
rect 354128 258068 354180 258120
rect 580172 258068 580224 258120
rect 3424 255212 3476 255264
rect 229468 255212 229520 255264
rect 3516 251132 3568 251184
rect 230388 251132 230440 251184
rect 353300 251132 353352 251184
rect 360844 251132 360896 251184
rect 353300 248344 353352 248396
rect 367744 248344 367796 248396
rect 32404 246984 32456 247036
rect 229836 246984 229888 247036
rect 385684 244264 385736 244316
rect 580172 244264 580224 244316
rect 353300 244196 353352 244248
rect 374644 244196 374696 244248
rect 22744 242836 22796 242888
rect 229652 242836 229704 242888
rect 353300 241408 353352 241460
rect 381544 241408 381596 241460
rect 14464 240048 14516 240100
rect 230388 240048 230440 240100
rect 353300 237328 353352 237380
rect 580356 237328 580408 237380
rect 7564 235900 7616 235952
rect 229836 235900 229888 235952
rect 353300 233180 353352 233232
rect 580448 233180 580500 233232
rect 3608 231752 3660 231804
rect 230388 231752 230440 231804
rect 353300 230392 353352 230444
rect 359464 230392 359516 230444
rect 3700 227672 3752 227724
rect 230388 227672 230440 227724
rect 353300 226244 353352 226296
rect 364984 226244 365036 226296
rect 43444 224884 43496 224936
rect 230388 224884 230440 224936
rect 353300 223524 353352 223576
rect 373264 223524 373316 223576
rect 25504 220736 25556 220788
rect 230388 220736 230440 220788
rect 353300 219308 353352 219360
rect 356704 219308 356756 219360
rect 353944 218016 353996 218068
rect 580172 218016 580224 218068
rect 17224 216588 17276 216640
rect 230388 216588 230440 216640
rect 353300 216588 353352 216640
rect 580448 216588 580500 216640
rect 8944 212440 8996 212492
rect 230388 212440 230440 212492
rect 353300 212440 353352 212492
rect 580632 212440 580684 212492
rect 3792 209720 3844 209772
rect 230020 209720 230072 209772
rect 353300 209312 353352 209364
rect 355324 209312 355376 209364
rect 3884 205572 3936 205624
rect 230388 205572 230440 205624
rect 353300 205572 353352 205624
rect 371884 205572 371936 205624
rect 31024 201424 31076 201476
rect 229652 201424 229704 201476
rect 353300 201424 353352 201476
rect 378784 201424 378836 201476
rect 353300 198636 353352 198688
rect 363604 198636 363656 198688
rect 26884 197276 26936 197328
rect 230388 197276 230440 197328
rect 18604 194488 18656 194540
rect 229652 194488 229704 194540
rect 353300 194488 353352 194540
rect 580724 194488 580776 194540
rect 10324 190408 10376 190460
rect 230388 190408 230440 190460
rect 353300 187620 353352 187672
rect 580816 187620 580868 187672
rect 3976 186260 4028 186312
rect 230388 186260 230440 186312
rect 353300 183472 353352 183524
rect 369124 183472 369176 183524
rect 4068 182112 4120 182164
rect 230388 182112 230440 182164
rect 353300 180752 353352 180804
rect 377404 180752 377456 180804
rect 221464 179324 221516 179376
rect 229652 179324 229704 179376
rect 354036 178032 354088 178084
rect 580172 178032 580224 178084
rect 353300 176604 353352 176656
rect 442264 176604 442316 176656
rect 28264 175176 28316 175228
rect 230388 175176 230440 175228
rect 353300 173816 353352 173868
rect 580908 173816 580960 173868
rect 21364 171028 21416 171080
rect 230388 171028 230440 171080
rect 13084 166948 13136 167000
rect 230388 166948 230440 167000
rect 353300 166948 353352 167000
rect 385684 166948 385736 167000
rect 3332 164160 3384 164212
rect 229652 164160 229704 164212
rect 353300 162800 353352 162852
rect 580264 162800 580316 162852
rect 3424 160012 3476 160064
rect 229468 160012 229520 160064
rect 3516 155864 3568 155916
rect 230388 155864 230440 155916
rect 353300 155864 353352 155916
rect 580356 155864 580408 155916
rect 353944 151784 353996 151836
rect 580172 151784 580224 151836
rect 3608 151716 3660 151768
rect 230388 151716 230440 151768
rect 353300 151716 353352 151768
rect 580448 151716 580500 151768
rect 3700 147568 3752 147620
rect 229652 147568 229704 147620
rect 3792 144848 3844 144900
rect 230388 144848 230440 144900
rect 353300 144848 353352 144900
rect 580540 144848 580592 144900
rect 3424 140700 3476 140752
rect 230388 140700 230440 140752
rect 353300 137980 353352 138032
rect 580172 137980 580224 138032
rect 3424 136552 3476 136604
rect 229836 136552 229888 136604
rect 3608 128324 3660 128376
rect 230388 128324 230440 128376
rect 354312 126896 354364 126948
rect 580172 126896 580224 126948
rect 3516 115948 3568 116000
rect 230204 115948 230256 116000
rect 353944 113092 353996 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 229744 111732 229796 111784
rect 3424 104864 3476 104916
rect 230388 104864 230440 104916
rect 354588 100648 354640 100700
rect 580172 100648 580224 100700
rect 238760 100104 238812 100156
rect 239220 100104 239272 100156
rect 285680 100104 285732 100156
rect 285956 100104 286008 100156
rect 225604 97928 225656 97980
rect 276848 97928 276900 97980
rect 284944 97928 284996 97980
rect 288808 97928 288860 97980
rect 334532 97928 334584 97980
rect 336188 97928 336240 97980
rect 257160 97860 257212 97912
rect 258632 97860 258684 97912
rect 268292 97792 268344 97844
rect 281264 97792 281316 97844
rect 341800 97792 341852 97844
rect 352564 97792 352616 97844
rect 224316 97724 224368 97776
rect 241060 97724 241112 97776
rect 255964 97724 256016 97776
rect 259368 97724 259420 97776
rect 275376 97724 275428 97776
rect 279332 97724 279384 97776
rect 322112 97724 322164 97776
rect 335636 97724 335688 97776
rect 349160 97724 349212 97776
rect 364984 97724 365036 97776
rect 221464 97656 221516 97708
rect 242532 97656 242584 97708
rect 345480 97656 345532 97708
rect 363604 97656 363656 97708
rect 224224 97588 224276 97640
rect 260288 97588 260340 97640
rect 228364 97520 228416 97572
rect 266636 97588 266688 97640
rect 274364 97588 274416 97640
rect 281724 97588 281776 97640
rect 294420 97588 294472 97640
rect 302240 97588 302292 97640
rect 317052 97588 317104 97640
rect 333336 97588 333388 97640
rect 335912 97588 335964 97640
rect 355324 97588 355376 97640
rect 275284 97520 275336 97572
rect 283472 97520 283524 97572
rect 295616 97520 295668 97572
rect 307208 97520 307260 97572
rect 311900 97520 311952 97572
rect 332140 97520 332192 97572
rect 338212 97520 338264 97572
rect 360844 97520 360896 97572
rect 295340 97452 295392 97504
rect 307024 97452 307076 97504
rect 330852 97452 330904 97504
rect 355508 97452 355560 97504
rect 124220 97384 124272 97436
rect 257620 97384 257672 97436
rect 276664 97384 276716 97436
rect 278044 97384 278096 97436
rect 279424 97384 279476 97436
rect 288532 97384 288584 97436
rect 297272 97384 297324 97436
rect 311164 97384 311216 97436
rect 331588 97384 331640 97436
rect 356704 97384 356756 97436
rect 106280 97316 106332 97368
rect 254032 97316 254084 97368
rect 269764 97316 269816 97368
rect 280804 97316 280856 97368
rect 300952 97316 301004 97368
rect 331864 97316 331916 97368
rect 335268 97316 335320 97368
rect 359464 97316 359516 97368
rect 10324 97248 10376 97300
rect 233056 97248 233108 97300
rect 257344 97248 257396 97300
rect 265164 97248 265216 97300
rect 298744 97248 298796 97300
rect 319444 97248 319496 97300
rect 332324 97248 332376 97300
rect 485044 97248 485096 97300
rect 303712 97180 303764 97232
rect 304448 97180 304500 97232
rect 350816 97112 350868 97164
rect 355416 97112 355468 97164
rect 242992 97044 243044 97096
rect 244740 97044 244792 97096
rect 279148 97044 279200 97096
rect 279884 97044 279936 97096
rect 295432 97044 295484 97096
rect 295892 97044 295944 97096
rect 296904 97044 296956 97096
rect 297364 97044 297416 97096
rect 301044 97044 301096 97096
rect 301504 97044 301556 97096
rect 303712 97044 303764 97096
rect 304172 97044 304224 97096
rect 305184 97044 305236 97096
rect 305644 97044 305696 97096
rect 327080 97044 327132 97096
rect 327540 97044 327592 97096
rect 328552 97044 328604 97096
rect 329012 97044 329064 97096
rect 231124 96976 231176 97028
rect 233516 96976 233568 97028
rect 233884 96976 233936 97028
rect 236460 96976 236512 97028
rect 278044 96976 278096 97028
rect 280528 96976 280580 97028
rect 298284 96976 298336 97028
rect 305736 96976 305788 97028
rect 325792 96976 325844 97028
rect 327724 96976 327776 97028
rect 328736 96976 328788 97028
rect 333244 96976 333296 97028
rect 348424 96976 348476 97028
rect 352748 96976 352800 97028
rect 231952 96908 232004 96960
rect 232780 96908 232832 96960
rect 233608 96908 233660 96960
rect 234252 96908 234304 96960
rect 234620 96908 234672 96960
rect 235356 96908 235408 96960
rect 237748 96908 237800 96960
rect 238024 96908 238076 96960
rect 239404 96908 239456 96960
rect 240324 96908 240376 96960
rect 242164 96908 242216 96960
rect 245476 96908 245528 96960
rect 255780 96908 255832 96960
rect 256148 96908 256200 96960
rect 256976 96908 257028 96960
rect 257252 96908 257304 96960
rect 259920 96908 259972 96960
rect 260380 96908 260432 96960
rect 261116 96908 261168 96960
rect 261392 96908 261444 96960
rect 262588 96908 262640 96960
rect 263324 96908 263376 96960
rect 275468 96908 275520 96960
rect 276112 96908 276164 96960
rect 276204 96908 276256 96960
rect 277308 96908 277360 96960
rect 279608 96908 279660 96960
rect 279884 96908 279936 96960
rect 281816 96908 281868 96960
rect 282184 96908 282236 96960
rect 283288 96908 283340 96960
rect 284024 96908 284076 96960
rect 284668 96908 284720 96960
rect 285220 96908 285272 96960
rect 286416 96908 286468 96960
rect 286692 96908 286744 96960
rect 287152 96908 287204 96960
rect 287428 96908 287480 96960
rect 287888 96908 287940 96960
rect 288164 96908 288216 96960
rect 290096 96908 290148 96960
rect 290832 96908 290884 96960
rect 291568 96908 291620 96960
rect 292396 96908 292448 96960
rect 292764 96908 292816 96960
rect 293132 96908 293184 96960
rect 294236 96908 294288 96960
rect 294696 96908 294748 96960
rect 295892 96908 295944 96960
rect 296536 96908 296588 96960
rect 297364 96908 297416 96960
rect 298008 96908 298060 96960
rect 298376 96908 298428 96960
rect 298836 96908 298888 96960
rect 299572 96908 299624 96960
rect 299940 96908 299992 96960
rect 300032 96908 300084 96960
rect 300676 96908 300728 96960
rect 302516 96908 302568 96960
rect 302976 96908 303028 96960
rect 304172 96908 304224 96960
rect 304816 96908 304868 96960
rect 305644 96908 305696 96960
rect 306288 96908 306340 96960
rect 306656 96908 306708 96960
rect 307484 96908 307536 96960
rect 307852 96908 307904 96960
rect 308588 96908 308640 96960
rect 309324 96908 309376 96960
rect 310060 96908 310112 96960
rect 310520 96908 310572 96960
rect 310888 96908 310940 96960
rect 312452 96908 312504 96960
rect 312728 96908 312780 96960
rect 313464 96908 313516 96960
rect 313832 96908 313884 96960
rect 313924 96908 313976 96960
rect 314200 96908 314252 96960
rect 314660 96908 314712 96960
rect 315764 96908 315816 96960
rect 316132 96908 316184 96960
rect 316592 96908 316644 96960
rect 317604 96908 317656 96960
rect 318524 96908 318576 96960
rect 318800 96908 318852 96960
rect 319536 96908 319588 96960
rect 321744 96908 321796 96960
rect 322572 96908 322624 96960
rect 322940 96908 322992 96960
rect 323308 96908 323360 96960
rect 323400 96908 323452 96960
rect 324044 96908 324096 96960
rect 324412 96908 324464 96960
rect 325516 96908 325568 96960
rect 327540 96908 327592 96960
rect 328184 96908 328236 96960
rect 329012 96908 329064 96960
rect 329656 96908 329708 96960
rect 330208 96908 330260 96960
rect 330484 96908 330536 96960
rect 332692 96908 332744 96960
rect 333520 96908 333572 96960
rect 334348 96908 334400 96960
rect 334992 96908 335044 96960
rect 335360 96908 335412 96960
rect 336464 96908 336516 96960
rect 337292 96908 337344 96960
rect 337660 96908 337712 96960
rect 338764 96908 338816 96960
rect 339224 96908 339276 96960
rect 339500 96908 339552 96960
rect 339868 96908 339920 96960
rect 339960 96908 340012 96960
rect 340604 96908 340656 96960
rect 341156 96908 341208 96960
rect 341432 96908 341484 96960
rect 342628 96908 342680 96960
rect 343364 96908 343416 96960
rect 344100 96908 344152 96960
rect 344744 96908 344796 96960
rect 345296 96908 345348 96960
rect 345940 96908 345992 96960
rect 346768 96908 346820 96960
rect 347412 96908 347464 96960
rect 347780 96908 347832 96960
rect 348608 96908 348660 96960
rect 349712 96908 349764 96960
rect 350172 96908 350224 96960
rect 350908 96908 350960 96960
rect 351184 96908 351236 96960
rect 235264 96840 235316 96892
rect 236736 96840 236788 96892
rect 240140 96840 240192 96892
rect 241428 96840 241480 96892
rect 243360 96840 243412 96892
rect 243728 96840 243780 96892
rect 255504 96840 255556 96892
rect 256240 96840 256292 96892
rect 260104 96840 260156 96892
rect 261024 96840 261076 96892
rect 261484 96840 261536 96892
rect 262956 96840 263008 96892
rect 270500 96840 270552 96892
rect 272524 96840 272576 96892
rect 275008 96840 275060 96892
rect 275744 96840 275796 96892
rect 279516 96840 279568 96892
rect 280252 96840 280304 96892
rect 287244 96840 287296 96892
rect 289084 96840 289136 96892
rect 290004 96840 290056 96892
rect 298100 96840 298152 96892
rect 299112 96840 299164 96892
rect 306380 96840 306432 96892
rect 307116 96840 307168 96892
rect 311992 96840 312044 96892
rect 313096 96840 313148 96892
rect 336832 96840 336884 96892
rect 337752 96840 337804 96892
rect 338488 96840 338540 96892
rect 339132 96840 339184 96892
rect 343640 96840 343692 96892
rect 344376 96840 344428 96892
rect 349436 96840 349488 96892
rect 350080 96840 350132 96892
rect 350632 96840 350684 96892
rect 352656 96840 352708 96892
rect 238024 96772 238076 96824
rect 238484 96772 238536 96824
rect 243544 96772 243596 96824
rect 244280 96772 244332 96824
rect 261392 96772 261444 96824
rect 261852 96772 261904 96824
rect 273996 96772 274048 96824
rect 274916 96772 274968 96824
rect 280804 96772 280856 96824
rect 284392 96772 284444 96824
rect 232504 96704 232556 96756
rect 234528 96704 234580 96756
rect 260196 96704 260248 96756
rect 262220 96704 262272 96756
rect 265440 96704 265492 96756
rect 267372 96704 267424 96756
rect 282184 96704 282236 96756
rect 283196 96704 283248 96756
rect 308220 96772 308272 96824
rect 315304 96772 315356 96824
rect 316316 96772 316368 96824
rect 323584 96772 323636 96824
rect 330116 96772 330168 96824
rect 332048 96772 332100 96824
rect 335636 96772 335688 96824
rect 336004 96772 336056 96824
rect 247684 96636 247736 96688
rect 248420 96636 248472 96688
rect 265624 96636 265676 96688
rect 268384 96636 268436 96688
rect 268476 96636 268528 96688
rect 271052 96636 271104 96688
rect 273904 96636 273956 96688
rect 274364 96636 274416 96688
rect 278136 96636 278188 96688
rect 281448 96636 281500 96688
rect 287244 96636 287296 96688
rect 340880 96636 340932 96688
rect 341892 96636 341944 96688
rect 209780 96160 209832 96212
rect 275192 96296 275244 96348
rect 201500 96092 201552 96144
rect 273720 96160 273772 96212
rect 307760 96160 307812 96212
rect 367100 96160 367152 96212
rect 308956 96092 309008 96144
rect 374000 96092 374052 96144
rect 182180 96024 182232 96076
rect 269580 96024 269632 96076
rect 321192 96024 321244 96076
rect 431960 96024 432012 96076
rect 80060 95956 80112 96008
rect 248604 95956 248656 96008
rect 333060 95956 333112 96008
rect 489920 95956 489972 96008
rect 4804 95888 4856 95940
rect 232136 95888 232188 95940
rect 300216 95888 300268 95940
rect 331220 95888 331272 95940
rect 344008 95888 344060 95940
rect 543740 95888 543792 95940
rect 326344 95752 326396 95804
rect 326804 95752 326856 95804
rect 257160 95412 257212 95464
rect 257344 95412 257396 95464
rect 284484 95344 284536 95396
rect 285588 95344 285640 95396
rect 310980 95344 311032 95396
rect 311256 95344 311308 95396
rect 268200 94800 268252 94852
rect 268660 94800 268712 94852
rect 264152 94732 264204 94784
rect 264520 94732 264572 94784
rect 267924 94732 267976 94784
rect 268568 94732 268620 94784
rect 305368 94732 305420 94784
rect 356060 94732 356112 94784
rect 227720 94664 227772 94716
rect 279056 94664 279108 94716
rect 306932 94664 306984 94716
rect 364340 94664 364392 94716
rect 195980 94596 196032 94648
rect 270500 94596 270552 94648
rect 311624 94596 311676 94648
rect 386420 94596 386472 94648
rect 125600 94528 125652 94580
rect 257896 94528 257948 94580
rect 263968 94528 264020 94580
rect 264520 94528 264572 94580
rect 266728 94528 266780 94580
rect 267096 94528 267148 94580
rect 269120 94528 269172 94580
rect 270132 94528 270184 94580
rect 270868 94528 270920 94580
rect 271604 94528 271656 94580
rect 272064 94528 272116 94580
rect 272708 94528 272760 94580
rect 333796 94528 333848 94580
rect 494060 94528 494112 94580
rect 60740 94460 60792 94512
rect 242992 94460 243044 94512
rect 246304 94460 246356 94512
rect 246672 94460 246724 94512
rect 247500 94460 247552 94512
rect 247960 94460 248012 94512
rect 248696 94460 248748 94512
rect 248972 94460 249024 94512
rect 250168 94460 250220 94512
rect 250444 94460 250496 94512
rect 251364 94460 251416 94512
rect 252100 94460 252152 94512
rect 252560 94460 252612 94512
rect 252836 94460 252888 94512
rect 267832 94460 267884 94512
rect 268660 94460 268712 94512
rect 270592 94460 270644 94512
rect 271328 94460 271380 94512
rect 346952 94460 347004 94512
rect 557540 94460 557592 94512
rect 247224 94392 247276 94444
rect 247868 94392 247920 94444
rect 248972 94324 249024 94376
rect 249432 94324 249484 94376
rect 250444 94324 250496 94376
rect 250904 94324 250956 94376
rect 270592 94324 270644 94376
rect 271512 94324 271564 94376
rect 304632 93372 304684 93424
rect 351920 93372 351972 93424
rect 200120 93304 200172 93356
rect 273260 93304 273312 93356
rect 332140 93304 332192 93356
rect 387800 93304 387852 93356
rect 193220 93236 193272 93288
rect 271972 93236 272024 93288
rect 326528 93236 326580 93288
rect 458180 93236 458232 93288
rect 160100 93168 160152 93220
rect 257436 93168 257488 93220
rect 336188 93168 336240 93220
rect 498200 93168 498252 93220
rect 71780 93100 71832 93152
rect 246764 93100 246816 93152
rect 351092 93100 351144 93152
rect 578240 93100 578292 93152
rect 215300 92012 215352 92064
rect 276388 92012 276440 92064
rect 207020 91944 207072 91996
rect 274640 91944 274692 91996
rect 305920 91944 305972 91996
rect 358820 91944 358872 91996
rect 164240 91876 164292 91928
rect 265900 91876 265952 91928
rect 312636 91876 312688 91928
rect 390560 91876 390612 91928
rect 113180 91808 113232 91860
rect 255412 91808 255464 91860
rect 336740 91808 336792 91860
rect 507860 91808 507912 91860
rect 46940 91740 46992 91792
rect 241888 91740 241940 91792
rect 344284 91740 344336 91792
rect 545120 91740 545172 91792
rect 213920 90516 213972 90568
rect 275468 90516 275520 90568
rect 306840 90516 306892 90568
rect 362960 90516 363012 90568
rect 171140 90448 171192 90500
rect 265440 90448 265492 90500
rect 313372 90448 313424 90500
rect 394700 90448 394752 90500
rect 151820 90380 151872 90432
rect 263048 90380 263100 90432
rect 337476 90380 337528 90432
rect 512000 90380 512052 90432
rect 26240 90312 26292 90364
rect 237472 90312 237524 90364
rect 347964 90312 348016 90364
rect 563060 90312 563112 90364
rect 265164 90108 265216 90160
rect 265532 90108 265584 90160
rect 220820 89156 220872 89208
rect 277676 89156 277728 89208
rect 315304 89156 315356 89208
rect 369860 89156 369912 89208
rect 175280 89088 175332 89140
rect 268108 89088 268160 89140
rect 319168 89088 319220 89140
rect 423680 89088 423732 89140
rect 147680 89020 147732 89072
rect 262496 89020 262548 89072
rect 325148 89020 325200 89072
rect 452660 89020 452712 89072
rect 16580 88952 16632 89004
rect 234620 88952 234672 89004
rect 338948 88952 339000 89004
rect 518900 88952 518952 89004
rect 230480 87796 230532 87848
rect 279884 87796 279936 87848
rect 309692 87796 309744 87848
rect 376760 87796 376812 87848
rect 178040 87728 178092 87780
rect 268200 87728 268252 87780
rect 322664 87728 322716 87780
rect 440332 87728 440384 87780
rect 139400 87660 139452 87712
rect 260840 87660 260892 87712
rect 330392 87660 330444 87712
rect 477500 87660 477552 87712
rect 103520 87592 103572 87644
rect 253480 87592 253532 87644
rect 267740 87592 267792 87644
rect 287244 87592 287296 87644
rect 339684 87592 339736 87644
rect 523040 87592 523092 87644
rect 354496 86912 354548 86964
rect 580172 86912 580224 86964
rect 219440 86436 219492 86488
rect 276204 86436 276256 86488
rect 184940 86368 184992 86420
rect 270316 86368 270368 86420
rect 306656 86368 306708 86420
rect 365720 86368 365772 86420
rect 146300 86300 146352 86352
rect 260196 86300 260248 86352
rect 323584 86300 323636 86352
rect 408500 86300 408552 86352
rect 20720 86232 20772 86284
rect 233884 86232 233936 86284
rect 316500 86232 316552 86284
rect 409880 86232 409932 86284
rect 3332 85484 3384 85536
rect 230112 85484 230164 85536
rect 308036 85008 308088 85060
rect 368480 85008 368532 85060
rect 218060 84940 218112 84992
rect 276940 84940 276992 84992
rect 311072 84940 311124 84992
rect 383660 84940 383712 84992
rect 202880 84872 202932 84924
rect 273812 84872 273864 84924
rect 340236 84872 340288 84924
rect 525800 84872 525852 84924
rect 107660 84804 107712 84856
rect 254308 84804 254360 84856
rect 294604 84804 294656 84856
rect 303620 84804 303672 84856
rect 347780 84804 347832 84856
rect 565820 84804 565872 84856
rect 310060 83648 310112 83700
rect 380900 83648 380952 83700
rect 189080 83580 189132 83632
rect 268476 83580 268528 83632
rect 355508 83580 355560 83632
rect 480260 83580 480312 83632
rect 126980 83512 127032 83564
rect 258172 83512 258224 83564
rect 327724 83512 327776 83564
rect 455420 83512 455472 83564
rect 85580 83444 85632 83496
rect 249800 83444 249852 83496
rect 267832 83444 267884 83496
rect 287428 83444 287480 83496
rect 349528 83444 349580 83496
rect 571340 83444 571392 83496
rect 193312 82220 193364 82272
rect 270868 82220 270920 82272
rect 312084 82220 312136 82272
rect 389180 82220 389232 82272
rect 129740 82152 129792 82204
rect 258724 82152 258776 82204
rect 333336 82152 333388 82204
rect 412640 82152 412692 82204
rect 89720 82084 89772 82136
rect 250168 82084 250220 82136
rect 302332 82084 302384 82136
rect 340880 82084 340932 82136
rect 340972 82084 341024 82136
rect 529940 82084 529992 82136
rect 308312 80860 308364 80912
rect 371240 80860 371292 80912
rect 211160 80792 211212 80844
rect 275560 80792 275612 80844
rect 314016 80792 314068 80844
rect 398840 80792 398892 80844
rect 128360 80724 128412 80776
rect 257344 80724 257396 80776
rect 326620 80724 326672 80776
rect 459560 80724 459612 80776
rect 78680 80656 78732 80708
rect 247684 80656 247736 80708
rect 256792 80656 256844 80708
rect 284760 80656 284812 80708
rect 342444 80656 342496 80708
rect 536840 80656 536892 80708
rect 224960 79500 225012 79552
rect 278228 79500 278280 79552
rect 150440 79432 150492 79484
rect 261484 79432 261536 79484
rect 312452 79432 312504 79484
rect 391940 79432 391992 79484
rect 53840 79364 53892 79416
rect 243268 79364 243320 79416
rect 317696 79364 317748 79416
rect 415400 79364 415452 79416
rect 13820 79296 13872 79348
rect 234896 79296 234948 79348
rect 343180 79296 343232 79348
rect 539600 79296 539652 79348
rect 197360 78072 197412 78124
rect 272064 78072 272116 78124
rect 316592 78072 316644 78124
rect 414020 78072 414072 78124
rect 132500 78004 132552 78056
rect 255964 78004 256016 78056
rect 320548 78004 320600 78056
rect 430580 78004 430632 78056
rect 100760 77936 100812 77988
rect 252652 77936 252704 77988
rect 344100 77936 344152 77988
rect 547880 77936 547932 77988
rect 231860 76712 231912 76764
rect 279700 76712 279752 76764
rect 168380 76644 168432 76696
rect 266820 76644 266872 76696
rect 324320 76644 324372 76696
rect 448520 76644 448572 76696
rect 41420 76576 41472 76628
rect 240416 76576 240468 76628
rect 331956 76576 332008 76628
rect 485780 76576 485832 76628
rect 7564 76508 7616 76560
rect 232228 76508 232280 76560
rect 346032 76508 346084 76560
rect 554780 76508 554832 76560
rect 304448 75352 304500 75404
rect 347780 75352 347832 75404
rect 173900 75284 173952 75336
rect 268660 75284 268712 75336
rect 312268 75284 312320 75336
rect 390652 75284 390704 75336
rect 135260 75216 135312 75268
rect 260012 75216 260064 75268
rect 330484 75216 330536 75268
rect 481640 75216 481692 75268
rect 40040 75148 40092 75200
rect 239404 75148 239456 75200
rect 347504 75148 347556 75200
rect 561680 75148 561732 75200
rect 305460 73992 305512 74044
rect 357440 73992 357492 74044
rect 180800 73924 180852 73976
rect 269396 73924 269448 73976
rect 309784 73924 309836 73976
rect 378140 73924 378192 73976
rect 143540 73856 143592 73908
rect 261116 73856 261168 73908
rect 323032 73856 323084 73908
rect 441620 73856 441672 73908
rect 35900 73788 35952 73840
rect 239496 73788 239548 73840
rect 352748 73788 352800 73840
rect 564532 73788 564584 73840
rect 354404 73108 354456 73160
rect 580172 73108 580224 73160
rect 198740 72564 198792 72616
rect 272800 72564 272852 72616
rect 305644 72564 305696 72616
rect 360200 72564 360252 72616
rect 153200 72496 153252 72548
rect 263600 72496 263652 72548
rect 310980 72496 311032 72548
rect 385040 72496 385092 72548
rect 29000 72428 29052 72480
rect 237748 72428 237800 72480
rect 328828 72428 328880 72480
rect 470600 72428 470652 72480
rect 3332 71680 3384 71732
rect 230020 71680 230072 71732
rect 310612 71136 310664 71188
rect 382280 71136 382332 71188
rect 201592 71068 201644 71120
rect 273444 71068 273496 71120
rect 325884 71068 325936 71120
rect 456892 71068 456944 71120
rect 121460 71000 121512 71052
rect 257068 71000 257120 71052
rect 303804 71000 303856 71052
rect 349160 71000 349212 71052
rect 349804 71000 349856 71052
rect 571984 71000 572036 71052
rect 209872 69776 209924 69828
rect 275100 69776 275152 69828
rect 309140 69776 309192 69828
rect 374092 69776 374144 69828
rect 157340 69708 157392 69760
rect 264336 69708 264388 69760
rect 321560 69708 321612 69760
rect 434720 69708 434772 69760
rect 110420 69640 110472 69692
rect 254768 69640 254820 69692
rect 302608 69640 302660 69692
rect 342260 69640 342312 69692
rect 352656 69640 352708 69692
rect 575480 69640 575532 69692
rect 216680 68416 216732 68468
rect 276480 68416 276532 68468
rect 314752 68416 314804 68468
rect 401600 68416 401652 68468
rect 161480 68348 161532 68400
rect 265256 68348 265308 68400
rect 332048 68348 332100 68400
rect 476120 68348 476172 68400
rect 93860 68280 93912 68332
rect 251180 68280 251232 68332
rect 335636 68280 335688 68332
rect 503720 68280 503772 68332
rect 165620 66988 165672 67040
rect 266084 66988 266136 67040
rect 315396 66988 315448 67040
rect 405740 66988 405792 67040
rect 95240 66920 95292 66972
rect 251732 66920 251784 66972
rect 332600 66920 332652 66972
rect 488540 66920 488592 66972
rect 69020 66852 69072 66904
rect 246028 66852 246080 66904
rect 265072 66852 265124 66904
rect 286508 66852 286560 66904
rect 296720 66852 296772 66904
rect 314752 66852 314804 66904
rect 342352 66852 342404 66904
rect 535460 66852 535512 66904
rect 172520 65628 172572 65680
rect 267464 65628 267516 65680
rect 318340 65628 318392 65680
rect 419540 65628 419592 65680
rect 82820 65560 82872 65612
rect 248696 65560 248748 65612
rect 333980 65560 334032 65612
rect 495440 65560 495492 65612
rect 44180 65492 44232 65544
rect 241244 65492 241296 65544
rect 348056 65492 348108 65544
rect 563704 65492 563756 65544
rect 179420 64268 179472 64320
rect 270132 64268 270184 64320
rect 316040 64268 316092 64320
rect 407120 64268 407172 64320
rect 88340 64200 88392 64252
rect 250260 64200 250312 64252
rect 319536 64200 319588 64252
rect 426440 64200 426492 64252
rect 57980 64132 58032 64184
rect 243820 64132 243872 64184
rect 341248 64132 341300 64184
rect 531320 64132 531372 64184
rect 183560 62908 183612 62960
rect 269672 62908 269724 62960
rect 307852 62908 307904 62960
rect 372620 62908 372672 62960
rect 74540 62840 74592 62892
rect 247408 62840 247460 62892
rect 321008 62840 321060 62892
rect 433340 62840 433392 62892
rect 64880 62772 64932 62824
rect 242164 62772 242216 62824
rect 345572 62772 345624 62824
rect 552020 62772 552072 62824
rect 186320 61480 186372 61532
rect 271328 61480 271380 61532
rect 306472 61480 306524 61532
rect 361580 61480 361632 61532
rect 63500 61412 63552 61464
rect 245108 61412 245160 61464
rect 336004 61412 336056 61464
rect 437480 61412 437532 61464
rect 11060 61344 11112 61396
rect 232504 61344 232556 61396
rect 346400 61344 346452 61396
rect 556160 61344 556212 61396
rect 354312 60664 354364 60716
rect 580172 60664 580224 60716
rect 208400 60120 208452 60172
rect 273996 60120 274048 60172
rect 301136 60120 301188 60172
rect 335452 60120 335504 60172
rect 149060 60052 149112 60104
rect 262680 60052 262732 60104
rect 313556 60052 313608 60104
rect 396080 60052 396132 60104
rect 12440 59984 12492 60036
rect 234804 59984 234856 60036
rect 318892 59984 318944 60036
rect 422300 59984 422352 60036
rect 222200 58760 222252 58812
rect 277768 58760 277820 58812
rect 321836 58760 321888 58812
rect 436100 58760 436152 58812
rect 131120 58692 131172 58744
rect 259000 58692 259052 58744
rect 323492 58692 323544 58744
rect 444380 58692 444432 58744
rect 84200 58624 84252 58676
rect 249248 58624 249300 58676
rect 298468 58624 298520 58676
rect 323032 58624 323084 58676
rect 349252 58624 349304 58676
rect 569960 58624 570012 58676
rect 314936 57332 314988 57384
rect 402980 57332 403032 57384
rect 133880 57264 133932 57316
rect 259644 57264 259696 57316
rect 324872 57264 324924 57316
rect 451280 57264 451332 57316
rect 73160 57196 73212 57248
rect 247040 57196 247092 57248
rect 338580 57196 338632 57248
rect 517520 57196 517572 57248
rect 317880 55972 317932 56024
rect 416780 55972 416832 56024
rect 143632 55904 143684 55956
rect 261668 55904 261720 55956
rect 327172 55904 327224 55956
rect 462320 55904 462372 55956
rect 62120 55836 62172 55888
rect 244832 55836 244884 55888
rect 343732 55836 343784 55888
rect 542360 55836 542412 55888
rect 320180 54612 320232 54664
rect 427820 54612 427872 54664
rect 127072 54544 127124 54596
rect 258448 54544 258500 54596
rect 327816 54544 327868 54596
rect 465172 54544 465224 54596
rect 77300 54476 77352 54528
rect 247224 54476 247276 54528
rect 349712 54476 349764 54528
rect 574100 54476 574152 54528
rect 162860 53116 162912 53168
rect 265164 53116 265216 53168
rect 324504 53116 324556 53168
rect 448612 53116 448664 53168
rect 114560 53048 114612 53100
rect 255596 53048 255648 53100
rect 300308 53048 300360 53100
rect 332600 53048 332652 53100
rect 333244 53048 333296 53100
rect 469220 53048 469272 53100
rect 167000 51756 167052 51808
rect 266452 51756 266504 51808
rect 322204 51756 322256 51808
rect 438860 51756 438912 51808
rect 8300 51688 8352 51740
rect 233700 51688 233752 51740
rect 329288 51688 329340 51740
rect 473360 51688 473412 51740
rect 169760 50396 169812 50448
rect 266728 50396 266780 50448
rect 323676 50396 323728 50448
rect 445760 50396 445812 50448
rect 66260 50328 66312 50380
rect 245752 50328 245804 50380
rect 331680 50328 331732 50380
rect 484400 50328 484452 50380
rect 229100 49104 229152 49156
rect 275376 49104 275428 49156
rect 111800 49036 111852 49088
rect 255044 49036 255096 49088
rect 331312 49036 331364 49088
rect 481732 49036 481784 49088
rect 2780 48968 2832 49020
rect 232596 48968 232648 49020
rect 333152 48968 333204 49020
rect 491300 48968 491352 49020
rect 176660 47608 176712 47660
rect 267924 47608 267976 47660
rect 334624 47608 334676 47660
rect 498292 47608 498344 47660
rect 59360 47540 59412 47592
rect 243544 47540 243596 47592
rect 337108 47540 337160 47592
rect 510620 47540 510672 47592
rect 354220 46860 354272 46912
rect 580172 46860 580224 46912
rect 187700 46316 187752 46368
rect 270684 46316 270736 46368
rect 99380 46248 99432 46300
rect 252836 46248 252888 46300
rect 303988 46248 304040 46300
rect 349252 46248 349304 46300
rect 33140 46180 33192 46232
rect 238852 46180 238904 46232
rect 334348 46180 334400 46232
rect 499580 46180 499632 46232
rect 3516 45500 3568 45552
rect 229928 45500 229980 45552
rect 226340 44888 226392 44940
rect 278872 44888 278924 44940
rect 335544 44888 335596 44940
rect 502340 44888 502392 44940
rect 60832 44820 60884 44872
rect 244556 44820 244608 44872
rect 338764 44820 338816 44872
rect 521660 44820 521712 44872
rect 191840 43460 191892 43512
rect 270592 43460 270644 43512
rect 335820 43460 335872 43512
rect 506480 43460 506532 43512
rect 48320 43392 48372 43444
rect 241980 43392 242032 43444
rect 340052 43392 340104 43444
rect 524420 43392 524472 43444
rect 194600 42168 194652 42220
rect 272156 42168 272208 42220
rect 110512 42100 110564 42152
rect 254584 42100 254636 42152
rect 336924 42100 336976 42152
rect 509240 42100 509292 42152
rect 52460 42032 52512 42084
rect 242624 42032 242676 42084
rect 301320 42032 301372 42084
rect 336740 42032 336792 42084
rect 341892 42032 341944 42084
rect 528560 42032 528612 42084
rect 205640 40808 205692 40860
rect 274272 40808 274324 40860
rect 81440 40740 81492 40792
rect 248788 40740 248840 40792
rect 337292 40740 337344 40792
rect 513380 40740 513432 40792
rect 44272 40672 44324 40724
rect 224316 40672 224368 40724
rect 342904 40672 342956 40724
rect 539692 40672 539744 40724
rect 223580 39448 223632 39500
rect 276664 39448 276716 39500
rect 302792 39448 302844 39500
rect 343732 39448 343784 39500
rect 67640 39380 67692 39432
rect 245844 39380 245896 39432
rect 338304 39380 338356 39432
rect 516140 39380 516192 39432
rect 6920 39312 6972 39364
rect 231124 39312 231176 39364
rect 343640 39312 343692 39364
rect 546500 39312 546552 39364
rect 135352 37952 135404 38004
rect 259828 37952 259880 38004
rect 338488 37952 338540 38004
rect 520280 37952 520332 38004
rect 102140 37884 102192 37936
rect 253020 37884 253072 37936
rect 345112 37884 345164 37936
rect 549260 37884 549312 37936
rect 138020 36592 138072 36644
rect 259920 36592 259972 36644
rect 339960 36592 340012 36644
rect 527180 36592 527232 36644
rect 22100 36524 22152 36576
rect 235264 36524 235316 36576
rect 345296 36524 345348 36576
rect 553400 36524 553452 36576
rect 142160 35232 142212 35284
rect 261208 35232 261260 35284
rect 341432 35232 341484 35284
rect 534080 35232 534132 35284
rect 17960 35164 18012 35216
rect 235356 35164 235408 35216
rect 346584 35164 346636 35216
rect 556252 35164 556304 35216
rect 151912 33804 151964 33856
rect 262588 33804 262640 33856
rect 342720 33804 342772 33856
rect 538220 33804 538272 33856
rect 98000 33736 98052 33788
rect 251364 33736 251416 33788
rect 348240 33736 348292 33788
rect 567200 33736 567252 33788
rect 3516 33056 3568 33108
rect 229836 33056 229888 33108
rect 354128 33056 354180 33108
rect 580172 33056 580224 33108
rect 304172 32444 304224 32496
rect 353300 32444 353352 32496
rect 118700 32376 118752 32428
rect 256976 32376 257028 32428
rect 314200 32376 314252 32428
rect 400220 32376 400272 32428
rect 305000 31152 305052 31204
rect 354680 31152 354732 31204
rect 155960 31084 156012 31136
rect 263784 31084 263836 31136
rect 318064 31084 318116 31136
rect 418160 31084 418212 31136
rect 109040 31016 109092 31068
rect 254400 31016 254452 31068
rect 342628 31016 342680 31068
rect 540980 31016 541032 31068
rect 160192 29656 160244 29708
rect 264980 29656 265032 29708
rect 315120 29656 315172 29708
rect 404360 29656 404412 29708
rect 104900 29588 104952 29640
rect 253572 29588 253624 29640
rect 301780 29588 301832 29640
rect 340972 29588 341024 29640
rect 345020 29588 345072 29640
rect 547972 29588 548024 29640
rect 96620 28296 96672 28348
rect 251916 28296 251968 28348
rect 316132 28296 316184 28348
rect 411260 28296 411312 28348
rect 56600 28228 56652 28280
rect 243360 28228 243412 28280
rect 302976 28228 303028 28280
rect 346400 28228 346452 28280
rect 347044 28228 347096 28280
rect 558920 28228 558972 28280
rect 212540 27004 212592 27056
rect 275008 27004 275060 27056
rect 102232 26936 102284 26988
rect 253112 26936 253164 26988
rect 310520 26936 310572 26988
rect 382372 26936 382424 26988
rect 55220 26868 55272 26920
rect 243452 26868 243504 26920
rect 300032 26868 300084 26920
rect 332876 26868 332928 26920
rect 349436 26868 349488 26920
rect 572812 26868 572864 26920
rect 185032 25576 185084 25628
rect 269856 25576 269908 25628
rect 313924 25576 313976 25628
rect 398932 25576 398984 25628
rect 86960 25508 87012 25560
rect 249984 25508 250036 25560
rect 327356 25508 327408 25560
rect 463700 25508 463752 25560
rect 154580 24148 154632 24200
rect 264520 24148 264572 24200
rect 314660 24148 314712 24200
rect 407212 24148 407264 24200
rect 27620 24080 27672 24132
rect 237656 24080 237708 24132
rect 327540 24080 327592 24132
rect 466460 24080 466512 24132
rect 176752 22788 176804 22840
rect 265624 22788 265676 22840
rect 317604 22788 317656 22840
rect 420920 22788 420972 22840
rect 93952 22720 94004 22772
rect 251640 22720 251692 22772
rect 329012 22720 329064 22772
rect 473452 22720 473504 22772
rect 158720 21428 158772 21480
rect 264060 21428 264112 21480
rect 319260 21428 319312 21480
rect 423772 21428 423824 21480
rect 122840 21360 122892 21412
rect 257988 21360 258040 21412
rect 260932 21360 260984 21412
rect 285956 21360 286008 21412
rect 332784 21360 332836 21412
rect 490012 21360 490064 21412
rect 354036 20612 354088 20664
rect 579988 20612 580040 20664
rect 297640 20068 297692 20120
rect 318892 20068 318944 20120
rect 144920 20000 144972 20052
rect 261392 20000 261444 20052
rect 306380 20000 306432 20052
rect 365812 20000 365864 20052
rect 30380 19932 30432 19984
rect 238300 19932 238352 19984
rect 258080 19932 258132 19984
rect 285036 19932 285088 19984
rect 318800 19932 318852 19984
rect 425060 19932 425112 19984
rect 118792 18640 118844 18692
rect 255504 18640 255556 18692
rect 320732 18640 320784 18692
rect 432052 18640 432104 18692
rect 49700 18572 49752 18624
rect 242256 18572 242308 18624
rect 242992 18572 243044 18624
rect 281816 18572 281868 18624
rect 296996 18572 297048 18624
rect 316040 18572 316092 18624
rect 332692 18572 332744 18624
rect 492680 18572 492732 18624
rect 226432 17348 226484 17400
rect 278412 17348 278464 17400
rect 85672 17280 85724 17332
rect 248972 17280 249024 17332
rect 311992 17280 312044 17332
rect 393320 17280 393372 17332
rect 2872 17212 2924 17264
rect 231952 17212 232004 17264
rect 301504 17212 301556 17264
rect 339592 17212 339644 17264
rect 355416 17212 355468 17264
rect 576860 17212 576912 17264
rect 205088 15920 205140 15972
rect 274088 15920 274140 15972
rect 339500 15920 339552 15972
rect 523776 15920 523828 15972
rect 69848 15852 69900 15904
rect 246396 15852 246448 15904
rect 299664 15852 299716 15904
rect 328736 15852 328788 15904
rect 346768 15852 346820 15904
rect 560392 15852 560444 15904
rect 298376 14560 298428 14612
rect 324596 14560 324648 14612
rect 116400 14492 116452 14544
rect 255872 14492 255924 14544
rect 277952 14492 278004 14544
rect 289176 14492 289228 14544
rect 317420 14492 317472 14544
rect 415492 14492 415544 14544
rect 53288 14424 53340 14476
rect 242900 14424 242952 14476
rect 251180 14424 251232 14476
rect 283564 14424 283616 14476
rect 305184 14424 305236 14476
rect 357532 14424 357584 14476
rect 364984 14424 365036 14476
rect 568672 14424 568724 14476
rect 270776 13200 270828 13252
rect 287704 13200 287756 13252
rect 309416 13200 309468 13252
rect 376024 13200 376076 13252
rect 190460 13132 190512 13184
rect 271236 13132 271288 13184
rect 320272 13132 320324 13184
rect 429200 13132 429252 13184
rect 91560 13064 91612 13116
rect 250720 13064 250772 13116
rect 252376 13064 252428 13116
rect 283840 13064 283892 13116
rect 302516 13064 302568 13116
rect 345296 13064 345348 13116
rect 363604 13064 363656 13116
rect 551008 13064 551060 13116
rect 75920 11772 75972 11824
rect 247592 11772 247644 11824
rect 264152 11772 264204 11824
rect 286232 11772 286284 11824
rect 309324 11772 309376 11824
rect 379520 11772 379572 11824
rect 71504 11704 71556 11756
rect 246304 11704 246356 11756
rect 247408 11704 247460 11756
rect 283012 11704 283064 11756
rect 301044 11704 301096 11756
rect 338672 11704 338724 11756
rect 352564 11704 352616 11756
rect 533712 11704 533764 11756
rect 160100 11636 160152 11688
rect 161296 11636 161348 11688
rect 176660 11636 176712 11688
rect 177856 11636 177908 11688
rect 184940 11636 184992 11688
rect 186136 11636 186188 11688
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 226340 11636 226392 11688
rect 227536 11636 227588 11688
rect 259460 10412 259512 10464
rect 284484 10412 284536 10464
rect 141240 10344 141292 10396
rect 260104 10344 260156 10396
rect 294696 10344 294748 10396
rect 306380 10344 306432 10396
rect 360844 10344 360896 10396
rect 515496 10344 515548 10396
rect 9680 10276 9732 10328
rect 233976 10276 234028 10328
rect 234620 10276 234672 10328
rect 279516 10276 279568 10328
rect 305736 10276 305788 10328
rect 321652 10276 321704 10328
rect 341156 10276 341208 10328
rect 532056 10276 532108 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 254676 9052 254728 9104
rect 280804 9052 280856 9104
rect 293776 9052 293828 9104
rect 300768 9052 300820 9104
rect 137652 8984 137704 9036
rect 224224 8984 224276 9036
rect 238116 8984 238168 9036
rect 280620 8984 280672 9036
rect 298100 8984 298152 9036
rect 326804 8984 326856 9036
rect 355324 8984 355376 9036
rect 505376 8984 505428 9036
rect 38384 8916 38436 8968
rect 239680 8916 239732 8968
rect 246396 8916 246448 8968
rect 282552 8916 282604 8968
rect 299480 8916 299532 8968
rect 328000 8916 328052 8968
rect 336832 8916 336884 8968
rect 514760 8916 514812 8968
rect 307116 8236 307168 8288
rect 309048 8236 309100 8288
rect 241704 7760 241756 7812
rect 273904 7760 273956 7812
rect 218152 7692 218204 7744
rect 225604 7692 225656 7744
rect 242900 7692 242952 7744
rect 281908 7692 281960 7744
rect 92756 7624 92808 7676
rect 250444 7624 250496 7676
rect 296168 7624 296220 7676
rect 312636 7624 312688 7676
rect 359464 7624 359516 7676
rect 501788 7624 501840 7676
rect 51356 7556 51408 7608
rect 221464 7556 221516 7608
rect 233424 7556 233476 7608
rect 279148 7556 279200 7608
rect 297364 7556 297416 7608
rect 320916 7556 320968 7608
rect 335360 7556 335412 7608
rect 507676 7556 507728 7608
rect 281908 6876 281960 6928
rect 289084 6876 289136 6928
rect 3424 6808 3476 6860
rect 229744 6808 229796 6860
rect 353944 6808 353996 6860
rect 580172 6808 580224 6860
rect 239312 6332 239364 6384
rect 268384 6332 268436 6384
rect 276020 6332 276072 6384
rect 284944 6332 284996 6384
rect 253480 6264 253532 6316
rect 283288 6264 283340 6316
rect 296904 6264 296956 6316
rect 318524 6264 318576 6316
rect 240508 6196 240560 6248
rect 278136 6196 278188 6248
rect 303712 6196 303764 6248
rect 351644 6196 351696 6248
rect 78588 6128 78640 6180
rect 247500 6128 247552 6180
rect 248788 6128 248840 6180
rect 282184 6128 282236 6180
rect 313464 6128 313516 6180
rect 397736 6128 397788 6180
rect 295892 6060 295944 6112
rect 313832 6060 313884 6112
rect 293500 5448 293552 5500
rect 299664 5448 299716 5500
rect 249984 4972 250036 5024
rect 275284 4972 275336 5024
rect 237012 4904 237064 4956
rect 269764 4904 269816 4956
rect 272432 4904 272484 4956
rect 287980 4904 288032 4956
rect 295708 4904 295760 4956
rect 310244 4904 310296 4956
rect 168472 4836 168524 4888
rect 228364 4836 228416 4888
rect 235816 4836 235868 4888
rect 278044 4836 278096 4888
rect 295432 4836 295484 4888
rect 311440 4836 311492 4888
rect 334164 4836 334216 4888
rect 34796 4768 34848 4820
rect 239220 4768 239272 4820
rect 245200 4768 245252 4820
rect 282276 4768 282328 4820
rect 299572 4768 299624 4820
rect 330392 4768 330444 4820
rect 356704 4836 356756 4888
rect 484032 4836 484084 4888
rect 497096 4768 497148 4820
rect 311164 4428 311216 4480
rect 317328 4428 317380 4480
rect 274824 4292 274876 4344
rect 279424 4292 279476 4344
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 193220 4156 193272 4208
rect 194416 4156 194468 4208
rect 218060 4156 218112 4208
rect 219256 4156 219308 4208
rect 307024 4156 307076 4208
rect 307944 4156 307996 4208
rect 319444 4156 319496 4208
rect 324320 4156 324372 4208
rect 331864 4156 331916 4208
rect 335084 4156 335136 4208
rect 485044 4156 485096 4208
rect 487620 4156 487672 4208
rect 43076 4088 43128 4140
rect 240692 4088 240744 4140
rect 284300 4088 284352 4140
rect 290372 4088 290424 4140
rect 292672 4088 292724 4140
rect 294880 4088 294932 4140
rect 324688 4088 324740 4140
rect 450912 4088 450964 4140
rect 39580 4020 39632 4072
rect 241428 4020 241480 4072
rect 283104 4020 283156 4072
rect 290188 4020 290240 4072
rect 292856 4020 292908 4072
rect 296076 4020 296128 4072
rect 324412 4020 324464 4072
rect 454500 4020 454552 4072
rect 35992 3952 36044 4004
rect 238760 3952 238812 4004
rect 292764 3952 292816 4004
rect 297272 3952 297324 4004
rect 326068 3952 326120 4004
rect 458088 3952 458140 4004
rect 32404 3884 32456 3936
rect 238024 3884 238076 3936
rect 279516 3884 279568 3936
rect 289360 3884 289412 3936
rect 293224 3884 293276 3936
rect 298468 3884 298520 3936
rect 326344 3884 326396 3936
rect 461584 3884 461636 3936
rect 28908 3816 28960 3868
rect 237840 3816 237892 3868
rect 277124 3816 277176 3868
rect 288624 3816 288676 3868
rect 293960 3816 294012 3868
rect 301964 3816 302016 3868
rect 327080 3816 327132 3868
rect 465172 3816 465224 3868
rect 25320 3748 25372 3800
rect 236920 3748 236972 3800
rect 273628 3748 273680 3800
rect 287888 3748 287940 3800
rect 328460 3748 328512 3800
rect 468668 3748 468720 3800
rect 24216 3680 24268 3732
rect 236828 3680 236880 3732
rect 267740 3680 267792 3732
rect 268476 3680 268528 3732
rect 270040 3680 270092 3732
rect 287152 3680 287204 3732
rect 328552 3680 328604 3732
rect 472256 3680 472308 3732
rect 572 3476 624 3528
rect 4804 3476 4856 3528
rect 5264 3476 5316 3528
rect 10324 3612 10376 3664
rect 19432 3612 19484 3664
rect 236000 3612 236052 3664
rect 266544 3612 266596 3664
rect 286416 3612 286468 3664
rect 329840 3612 329892 3664
rect 475752 3612 475804 3664
rect 7564 3544 7616 3596
rect 20628 3544 20680 3596
rect 236276 3544 236328 3596
rect 262956 3544 263008 3596
rect 285680 3544 285732 3596
rect 286600 3544 286652 3596
rect 290096 3544 290148 3596
rect 291568 3544 291620 3596
rect 293684 3544 293736 3596
rect 321744 3544 321796 3596
rect 1676 3272 1728 3324
rect 15936 3476 15988 3528
rect 235080 3476 235132 3528
rect 259460 3476 259512 3528
rect 260656 3476 260708 3528
rect 285404 3476 285456 3528
rect 290556 3476 290608 3528
rect 11152 3408 11204 3460
rect 233608 3408 233660 3460
rect 255872 3408 255924 3460
rect 285220 3408 285272 3460
rect 292028 3408 292080 3460
rect 292580 3408 292632 3460
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 46664 3340 46716 3392
rect 241520 3340 241572 3392
rect 259460 3340 259512 3392
rect 285312 3340 285364 3392
rect 294236 3340 294288 3392
rect 305552 3340 305604 3392
rect 60740 3272 60792 3324
rect 61660 3272 61712 3324
rect 85580 3272 85632 3324
rect 86500 3272 86552 3324
rect 110420 3272 110472 3324
rect 111616 3272 111668 3324
rect 118700 3272 118752 3324
rect 119896 3272 119948 3324
rect 117596 3204 117648 3256
rect 255780 3272 255832 3324
rect 280712 3272 280764 3324
rect 289636 3272 289688 3324
rect 290188 3272 290240 3324
rect 291660 3272 291712 3324
rect 121092 3204 121144 3256
rect 257252 3204 257304 3256
rect 351184 3544 351236 3596
rect 582196 3544 582248 3596
rect 330208 3476 330260 3528
rect 479340 3476 479392 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 563704 3476 563756 3528
rect 564440 3476 564492 3528
rect 571984 3476 572036 3528
rect 572720 3476 572772 3528
rect 349252 3408 349304 3460
rect 350448 3408 350500 3460
rect 350908 3408 350960 3460
rect 581000 3408 581052 3460
rect 323400 3340 323452 3392
rect 447416 3340 447468 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 322940 3272 322992 3324
rect 443828 3272 443880 3324
rect 440240 3204 440292 3256
rect 440332 3204 440384 3256
rect 441528 3204 441580 3256
rect 168380 3136 168432 3188
rect 169576 3136 169628 3188
rect 288992 3136 289044 3188
rect 291292 3136 291344 3188
rect 357532 3136 357584 3188
rect 358728 3136 358780 3188
rect 374092 3136 374144 3188
rect 375288 3136 375340 3188
rect 382372 3136 382424 3188
rect 383568 3136 383620 3188
rect 398932 3136 398984 3188
rect 400128 3136 400180 3188
rect 407120 3136 407172 3188
rect 408408 3136 408460 3188
rect 415400 3136 415452 3188
rect 416688 3136 416740 3188
rect 423772 3136 423824 3188
rect 424968 3136 425020 3188
rect 431960 3136 432012 3188
rect 433248 3136 433300 3188
rect 287796 3068 287848 3120
rect 291200 3068 291252 3120
rect 340880 2728 340932 2780
rect 342168 2728 342220 2780
rect 365720 1504 365772 1556
rect 367008 1504 367060 1556
rect 390560 1504 390612 1556
rect 391848 1504 391900 1556
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3332 632120 3384 632126
rect 3330 632088 3332 632097
rect 3384 632088 3386 632097
rect 3330 632023 3386 632032
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3344 618322 3372 619103
rect 3332 618316 3384 618322
rect 3332 618258 3384 618264
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3160 579834 3188 579935
rect 3148 579828 3200 579834
rect 3148 579770 3200 579776
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 475250 3372 475623
rect 3332 475244 3384 475250
rect 3332 475186 3384 475192
rect 2962 423600 3018 423609
rect 2962 423535 3018 423544
rect 2976 422346 3004 423535
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3160 318850 3188 319223
rect 3148 318844 3200 318850
rect 3148 318786 3200 318792
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3344 305046 3372 306167
rect 3332 305040 3384 305046
rect 3332 304982 3384 304988
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3252 266422 3280 267135
rect 3240 266416 3292 266422
rect 3240 266358 3292 266364
rect 3436 255270 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3344 164218 3372 254079
rect 3528 251190 3556 658135
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3516 251184 3568 251190
rect 3516 251126 3568 251132
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3436 160070 3464 241023
rect 3620 231810 3648 566879
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3608 231804 3660 231810
rect 3608 231746 3660 231752
rect 3712 227730 3740 553823
rect 3790 462632 3846 462641
rect 3790 462567 3846 462576
rect 3700 227724 3752 227730
rect 3700 227666 3752 227672
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 3424 160064 3476 160070
rect 3424 160006 3476 160012
rect 3528 155922 3556 214911
rect 3804 209778 3832 462567
rect 3882 449576 3938 449585
rect 3882 449511 3938 449520
rect 3792 209772 3844 209778
rect 3792 209714 3844 209720
rect 3896 205630 3924 449511
rect 3974 358456 4030 358465
rect 3974 358391 4030 358400
rect 3884 205624 3936 205630
rect 3884 205566 3936 205572
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3516 155916 3568 155922
rect 3516 155858 3568 155864
rect 3620 151774 3648 201855
rect 3698 188864 3754 188873
rect 3698 188799 3754 188808
rect 3608 151768 3660 151774
rect 3608 151710 3660 151716
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 140758 3464 149767
rect 3712 147626 3740 188799
rect 3988 186318 4016 358391
rect 4066 345400 4122 345409
rect 4066 345335 4122 345344
rect 3976 186312 4028 186318
rect 3976 186254 4028 186260
rect 4080 182170 4108 345335
rect 4816 259418 4844 683674
rect 6932 262886 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 22744 618316 22796 618322
rect 22744 618258 22796 618264
rect 14464 605872 14516 605878
rect 14464 605814 14516 605820
rect 7564 579828 7616 579834
rect 7564 579770 7616 579776
rect 6920 262880 6972 262886
rect 6920 262822 6972 262828
rect 4804 259412 4856 259418
rect 4804 259354 4856 259360
rect 7576 235958 7604 579770
rect 8944 475244 8996 475250
rect 8944 475186 8996 475192
rect 7564 235952 7616 235958
rect 7564 235894 7616 235900
rect 8956 212498 8984 475186
rect 10324 371272 10376 371278
rect 10324 371214 10376 371220
rect 8944 212492 8996 212498
rect 8944 212434 8996 212440
rect 10336 190466 10364 371214
rect 13084 266416 13136 266422
rect 13084 266358 13136 266364
rect 10324 190460 10376 190466
rect 10324 190402 10376 190408
rect 4068 182164 4120 182170
rect 4068 182106 4120 182112
rect 13096 167006 13124 266358
rect 14476 240106 14504 605814
rect 17224 501016 17276 501022
rect 17224 500958 17276 500964
rect 14464 240100 14516 240106
rect 14464 240042 14516 240048
rect 17236 216646 17264 500958
rect 18604 397520 18656 397526
rect 18604 397462 18656 397468
rect 17224 216640 17276 216646
rect 17224 216582 17276 216588
rect 18616 194546 18644 397462
rect 21364 292596 21416 292602
rect 21364 292538 21416 292544
rect 18604 194540 18656 194546
rect 18604 194482 18656 194488
rect 21376 171086 21404 292538
rect 22756 242894 22784 618258
rect 23492 262954 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 32404 632120 32456 632126
rect 32404 632062 32456 632068
rect 25504 514820 25556 514826
rect 25504 514762 25556 514768
rect 23480 262948 23532 262954
rect 23480 262890 23532 262896
rect 22744 242888 22796 242894
rect 22744 242830 22796 242836
rect 25516 220794 25544 514762
rect 31024 422340 31076 422346
rect 31024 422282 31076 422288
rect 26884 409896 26936 409902
rect 26884 409838 26936 409844
rect 25504 220788 25556 220794
rect 25504 220730 25556 220736
rect 26896 197334 26924 409838
rect 28264 305040 28316 305046
rect 28264 304982 28316 304988
rect 26884 197328 26936 197334
rect 26884 197270 26936 197276
rect 28276 175234 28304 304982
rect 31036 201482 31064 422282
rect 32416 247042 32444 632062
rect 40052 263022 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 43444 527196 43496 527202
rect 43444 527138 43496 527144
rect 40040 263016 40092 263022
rect 40040 262958 40092 262964
rect 32404 247036 32456 247042
rect 32404 246978 32456 246984
rect 43456 224942 43484 527138
rect 71792 263090 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 263158 88380 702406
rect 104912 263226 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 263294 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 263362 153240 702406
rect 169772 263430 169800 702406
rect 201512 263498 201540 702986
rect 218072 263566 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 221464 318844 221516 318850
rect 221464 318786 221516 318792
rect 218060 263560 218112 263566
rect 218060 263502 218112 263508
rect 201500 263492 201552 263498
rect 201500 263434 201552 263440
rect 169760 263424 169812 263430
rect 169760 263366 169812 263372
rect 153200 263356 153252 263362
rect 153200 263298 153252 263304
rect 136640 263288 136692 263294
rect 136640 263230 136692 263236
rect 104900 263220 104952 263226
rect 104900 263162 104952 263168
rect 88340 263152 88392 263158
rect 88340 263094 88392 263100
rect 71780 263084 71832 263090
rect 71780 263026 71832 263032
rect 43444 224936 43496 224942
rect 43444 224878 43496 224884
rect 31024 201476 31076 201482
rect 31024 201418 31076 201424
rect 221476 179382 221504 318786
rect 234632 262886 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700330 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 279424 700324 279476 700330
rect 279424 700266 279476 700272
rect 278596 263560 278648 263566
rect 278596 263502 278648 263508
rect 274180 263492 274232 263498
rect 274180 263434 274232 263440
rect 269764 263424 269816 263430
rect 269764 263366 269816 263372
rect 265348 263356 265400 263362
rect 265348 263298 265400 263304
rect 260840 263288 260892 263294
rect 260840 263230 260892 263236
rect 256424 263220 256476 263226
rect 256424 263162 256476 263168
rect 252008 263152 252060 263158
rect 252008 263094 252060 263100
rect 247500 263084 247552 263090
rect 247500 263026 247552 263032
rect 243084 263016 243136 263022
rect 243084 262958 243136 262964
rect 238668 262948 238720 262954
rect 238668 262890 238720 262896
rect 234252 262880 234304 262886
rect 234252 262822 234304 262828
rect 234620 262880 234672 262886
rect 234620 262822 234672 262828
rect 234264 259964 234292 262822
rect 238680 259964 238708 262890
rect 243096 259964 243124 262958
rect 247512 259964 247540 263026
rect 252020 259964 252048 263094
rect 256436 259964 256464 263162
rect 260852 259964 260880 263230
rect 265360 259964 265388 263298
rect 269776 259964 269804 263366
rect 274192 259964 274220 263434
rect 278608 259964 278636 263502
rect 279436 262954 279464 700266
rect 282932 263022 282960 702406
rect 300136 700330 300164 703520
rect 309140 700936 309192 700942
rect 309140 700878 309192 700884
rect 300860 700392 300912 700398
rect 300860 700334 300912 700340
rect 295340 700324 295392 700330
rect 295340 700266 295392 700272
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 295352 267734 295380 700266
rect 295352 267706 296024 267734
rect 282920 263016 282972 263022
rect 282920 262958 282972 262964
rect 291936 263016 291988 263022
rect 291936 262958 291988 262964
rect 279424 262948 279476 262954
rect 279424 262890 279476 262896
rect 287520 262948 287572 262954
rect 287520 262890 287572 262896
rect 283104 262880 283156 262886
rect 283104 262822 283156 262828
rect 283116 259964 283144 262822
rect 287532 259964 287560 262890
rect 291948 259964 291976 262958
rect 295996 259978 296024 267706
rect 295996 259950 296470 259978
rect 300872 259964 300900 700334
rect 305000 700324 305052 700330
rect 305000 700266 305052 700272
rect 305012 259978 305040 700266
rect 309152 267734 309180 700878
rect 313280 700868 313332 700874
rect 313280 700810 313332 700816
rect 313292 267734 313320 700810
rect 317420 700800 317472 700806
rect 317420 700742 317472 700748
rect 317432 267734 317460 700742
rect 322940 700732 322992 700738
rect 322940 700674 322992 700680
rect 322952 267734 322980 700674
rect 327080 700664 327132 700670
rect 327080 700606 327132 700612
rect 309152 267706 309456 267734
rect 313292 267706 313872 267734
rect 317432 267706 318288 267734
rect 322952 267706 323072 267734
rect 309428 259978 309456 267706
rect 313844 259978 313872 267706
rect 318260 259978 318288 267706
rect 305012 259950 305302 259978
rect 309428 259950 309810 259978
rect 313844 259950 314226 259978
rect 318260 259950 318642 259978
rect 323044 259964 323072 267706
rect 327092 259978 327120 700606
rect 331312 700596 331364 700602
rect 331312 700538 331364 700544
rect 331324 267734 331352 700538
rect 332520 700398 332548 703520
rect 335360 700528 335412 700534
rect 335360 700470 335412 700476
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 335372 267734 335400 700470
rect 340880 700460 340932 700466
rect 340880 700402 340932 700408
rect 331324 267706 331536 267734
rect 335372 267706 335952 267734
rect 331508 259978 331536 267706
rect 335924 259978 335952 267706
rect 327092 259950 327566 259978
rect 331508 259950 331982 259978
rect 335924 259950 336398 259978
rect 340892 259964 340920 700402
rect 345020 700392 345072 700398
rect 345020 700334 345072 700340
rect 345032 259978 345060 700334
rect 348804 700330 348832 703520
rect 364996 700942 365024 703520
rect 364984 700936 365036 700942
rect 364984 700878 365036 700884
rect 397472 700874 397500 703520
rect 397460 700868 397512 700874
rect 397460 700810 397512 700816
rect 413664 700806 413692 703520
rect 413652 700800 413704 700806
rect 413652 700742 413704 700748
rect 429856 700738 429884 703520
rect 429844 700732 429896 700738
rect 429844 700674 429896 700680
rect 462332 700670 462360 703520
rect 462320 700664 462372 700670
rect 462320 700606 462372 700612
rect 478524 700602 478552 703520
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 494808 700534 494836 703520
rect 494796 700528 494848 700534
rect 494796 700470 494848 700476
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700398 543504 703520
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 559668 700330 559696 703520
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 349160 700324 349212 700330
rect 349160 700266 349212 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 349172 267734 349200 700266
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 353944 683188 353996 683194
rect 353944 683130 353996 683136
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 349172 267706 349384 267734
rect 349356 259978 349384 267706
rect 345032 259950 345322 259978
rect 349356 259950 349738 259978
rect 229100 259412 229152 259418
rect 229100 259354 229152 259360
rect 229112 258097 229140 259354
rect 229098 258088 229154 258097
rect 229098 258023 229154 258032
rect 229468 255264 229520 255270
rect 229468 255206 229520 255212
rect 229480 254289 229508 255206
rect 353956 254561 353984 683130
rect 360844 670744 360896 670750
rect 580172 670744 580224 670750
rect 360844 670686 360896 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 359464 563100 359516 563106
rect 359464 563042 359516 563048
rect 356704 510672 356756 510678
rect 356704 510614 356756 510620
rect 355324 456816 355376 456822
rect 355324 456758 355376 456764
rect 354036 364404 354088 364410
rect 354036 364346 354088 364352
rect 353942 254552 353998 254561
rect 353942 254487 353998 254496
rect 229466 254280 229522 254289
rect 229466 254215 229522 254224
rect 230388 251184 230440 251190
rect 230388 251126 230440 251132
rect 353300 251184 353352 251190
rect 353300 251126 353352 251132
rect 230400 250481 230428 251126
rect 353312 251025 353340 251126
rect 353298 251016 353354 251025
rect 353298 250951 353354 250960
rect 230386 250472 230442 250481
rect 230386 250407 230442 250416
rect 353300 248396 353352 248402
rect 353300 248338 353352 248344
rect 353312 247489 353340 248338
rect 353298 247480 353354 247489
rect 353298 247415 353354 247424
rect 229836 247036 229888 247042
rect 229836 246978 229888 246984
rect 229848 246673 229876 246978
rect 229834 246664 229890 246673
rect 229834 246599 229890 246608
rect 353300 244248 353352 244254
rect 353300 244190 353352 244196
rect 353312 243953 353340 244190
rect 353298 243944 353354 243953
rect 353298 243879 353354 243888
rect 229652 242888 229704 242894
rect 229650 242856 229652 242865
rect 229704 242856 229706 242865
rect 229650 242791 229706 242800
rect 353300 241460 353352 241466
rect 353300 241402 353352 241408
rect 353312 240417 353340 241402
rect 353298 240408 353354 240417
rect 353298 240343 353354 240352
rect 230388 240100 230440 240106
rect 230388 240042 230440 240048
rect 230400 239057 230428 240042
rect 230386 239048 230442 239057
rect 230386 238983 230442 238992
rect 353300 237380 353352 237386
rect 353300 237322 353352 237328
rect 353312 236881 353340 237322
rect 353298 236872 353354 236881
rect 353298 236807 353354 236816
rect 229836 235952 229888 235958
rect 229836 235894 229888 235900
rect 229848 235249 229876 235894
rect 229834 235240 229890 235249
rect 229834 235175 229890 235184
rect 353300 233232 353352 233238
rect 353298 233200 353300 233209
rect 353352 233200 353354 233209
rect 353298 233135 353354 233144
rect 230388 231804 230440 231810
rect 230388 231746 230440 231752
rect 230400 231441 230428 231746
rect 230386 231432 230442 231441
rect 230386 231367 230442 231376
rect 353300 230444 353352 230450
rect 353300 230386 353352 230392
rect 353312 229673 353340 230386
rect 353298 229664 353354 229673
rect 353298 229599 353354 229608
rect 230388 227724 230440 227730
rect 230388 227666 230440 227672
rect 230400 227633 230428 227666
rect 230386 227624 230442 227633
rect 230386 227559 230442 227568
rect 353300 226296 353352 226302
rect 353300 226238 353352 226244
rect 353312 226137 353340 226238
rect 353298 226128 353354 226137
rect 353298 226063 353354 226072
rect 230388 224936 230440 224942
rect 230388 224878 230440 224884
rect 230400 223825 230428 224878
rect 230386 223816 230442 223825
rect 230386 223751 230442 223760
rect 353300 223576 353352 223582
rect 353300 223518 353352 223524
rect 353312 222601 353340 223518
rect 353298 222592 353354 222601
rect 353298 222527 353354 222536
rect 230388 220788 230440 220794
rect 230388 220730 230440 220736
rect 230400 220017 230428 220730
rect 230386 220008 230442 220017
rect 230386 219943 230442 219952
rect 353300 219360 353352 219366
rect 353300 219302 353352 219308
rect 353312 219065 353340 219302
rect 353298 219056 353354 219065
rect 353298 218991 353354 219000
rect 353944 218068 353996 218074
rect 353944 218010 353996 218016
rect 230388 216640 230440 216646
rect 230388 216582 230440 216588
rect 353300 216640 353352 216646
rect 353300 216582 353352 216588
rect 230400 216209 230428 216582
rect 230386 216200 230442 216209
rect 230386 216135 230442 216144
rect 353312 215529 353340 216582
rect 353298 215520 353354 215529
rect 353298 215455 353354 215464
rect 230388 212492 230440 212498
rect 230388 212434 230440 212440
rect 353300 212492 353352 212498
rect 353300 212434 353352 212440
rect 230400 212401 230428 212434
rect 230386 212392 230442 212401
rect 230386 212327 230442 212336
rect 353312 211993 353340 212434
rect 353298 211984 353354 211993
rect 353298 211919 353354 211928
rect 230020 209772 230072 209778
rect 230020 209714 230072 209720
rect 230032 208593 230060 209714
rect 353300 209364 353352 209370
rect 353300 209306 353352 209312
rect 230018 208584 230074 208593
rect 230018 208519 230074 208528
rect 353312 208457 353340 209306
rect 353298 208448 353354 208457
rect 353298 208383 353354 208392
rect 230388 205624 230440 205630
rect 230388 205566 230440 205572
rect 353300 205624 353352 205630
rect 353300 205566 353352 205572
rect 230400 204785 230428 205566
rect 353312 204785 353340 205566
rect 230386 204776 230442 204785
rect 230386 204711 230442 204720
rect 353298 204776 353354 204785
rect 353298 204711 353354 204720
rect 229652 201476 229704 201482
rect 229652 201418 229704 201424
rect 353300 201476 353352 201482
rect 353300 201418 353352 201424
rect 229664 200977 229692 201418
rect 353312 201249 353340 201418
rect 353298 201240 353354 201249
rect 353298 201175 353354 201184
rect 229650 200968 229706 200977
rect 229650 200903 229706 200912
rect 353300 198688 353352 198694
rect 353300 198630 353352 198636
rect 353312 197713 353340 198630
rect 353298 197704 353354 197713
rect 353298 197639 353354 197648
rect 230388 197328 230440 197334
rect 230388 197270 230440 197276
rect 230400 197169 230428 197270
rect 230386 197160 230442 197169
rect 230386 197095 230442 197104
rect 229652 194540 229704 194546
rect 229652 194482 229704 194488
rect 353300 194540 353352 194546
rect 353300 194482 353352 194488
rect 229664 193361 229692 194482
rect 353312 194177 353340 194482
rect 353298 194168 353354 194177
rect 353298 194103 353354 194112
rect 229650 193352 229706 193361
rect 229650 193287 229706 193296
rect 230388 190460 230440 190466
rect 230388 190402 230440 190408
rect 230400 189553 230428 190402
rect 230386 189544 230442 189553
rect 230386 189479 230442 189488
rect 353300 187672 353352 187678
rect 353300 187614 353352 187620
rect 353312 187105 353340 187614
rect 353298 187096 353354 187105
rect 353298 187031 353354 187040
rect 230388 186312 230440 186318
rect 230388 186254 230440 186260
rect 230400 185745 230428 186254
rect 230386 185736 230442 185745
rect 230386 185671 230442 185680
rect 353298 183560 353354 183569
rect 353298 183495 353300 183504
rect 353352 183495 353354 183504
rect 353300 183466 353352 183472
rect 230388 182164 230440 182170
rect 230388 182106 230440 182112
rect 230400 181937 230428 182106
rect 230386 181928 230442 181937
rect 230386 181863 230442 181872
rect 353300 180804 353352 180810
rect 353300 180746 353352 180752
rect 353312 179897 353340 180746
rect 353298 179888 353354 179897
rect 353298 179823 353354 179832
rect 221464 179376 221516 179382
rect 221464 179318 221516 179324
rect 229652 179376 229704 179382
rect 229652 179318 229704 179324
rect 229664 178129 229692 179318
rect 229650 178120 229706 178129
rect 229650 178055 229706 178064
rect 353300 176656 353352 176662
rect 353300 176598 353352 176604
rect 353312 176361 353340 176598
rect 353298 176352 353354 176361
rect 353298 176287 353354 176296
rect 28264 175228 28316 175234
rect 28264 175170 28316 175176
rect 230388 175228 230440 175234
rect 230388 175170 230440 175176
rect 230400 174321 230428 175170
rect 230386 174312 230442 174321
rect 230386 174247 230442 174256
rect 353300 173868 353352 173874
rect 353300 173810 353352 173816
rect 353312 172825 353340 173810
rect 353298 172816 353354 172825
rect 353298 172751 353354 172760
rect 21364 171080 21416 171086
rect 21364 171022 21416 171028
rect 230388 171080 230440 171086
rect 230388 171022 230440 171028
rect 230400 170513 230428 171022
rect 230386 170504 230442 170513
rect 230386 170439 230442 170448
rect 13084 167000 13136 167006
rect 13084 166942 13136 166948
rect 230388 167000 230440 167006
rect 230388 166942 230440 166948
rect 353300 167000 353352 167006
rect 353300 166942 353352 166948
rect 230400 166705 230428 166942
rect 230386 166696 230442 166705
rect 230386 166631 230442 166640
rect 353312 165753 353340 166942
rect 353298 165744 353354 165753
rect 353298 165679 353354 165688
rect 229652 164212 229704 164218
rect 229652 164154 229704 164160
rect 229664 162897 229692 164154
rect 3790 162888 3846 162897
rect 3790 162823 3846 162832
rect 229650 162888 229706 162897
rect 229650 162823 229706 162832
rect 353300 162852 353352 162858
rect 3700 147620 3752 147626
rect 3700 147562 3752 147568
rect 3804 144906 3832 162823
rect 353300 162794 353352 162800
rect 353312 162217 353340 162794
rect 353298 162208 353354 162217
rect 353298 162143 353354 162152
rect 229468 160064 229520 160070
rect 229468 160006 229520 160012
rect 229480 159089 229508 160006
rect 229466 159080 229522 159089
rect 229466 159015 229522 159024
rect 353956 158681 353984 218010
rect 354048 190641 354076 364346
rect 354312 259412 354364 259418
rect 354312 259354 354364 259360
rect 354324 258233 354352 259354
rect 354310 258224 354366 258233
rect 354310 258159 354366 258168
rect 354128 258120 354180 258126
rect 354128 258062 354180 258068
rect 354034 190632 354090 190641
rect 354034 190567 354090 190576
rect 354036 178084 354088 178090
rect 354036 178026 354088 178032
rect 353942 158672 353998 158681
rect 353942 158607 353998 158616
rect 230388 155916 230440 155922
rect 230388 155858 230440 155864
rect 353300 155916 353352 155922
rect 353300 155858 353352 155864
rect 230400 155281 230428 155858
rect 230386 155272 230442 155281
rect 230386 155207 230442 155216
rect 353312 155145 353340 155858
rect 353298 155136 353354 155145
rect 353298 155071 353354 155080
rect 353944 151836 353996 151842
rect 353944 151778 353996 151784
rect 230388 151768 230440 151774
rect 230388 151710 230440 151716
rect 353300 151768 353352 151774
rect 353300 151710 353352 151716
rect 230400 151473 230428 151710
rect 353312 151473 353340 151710
rect 230386 151464 230442 151473
rect 230386 151399 230442 151408
rect 353298 151464 353354 151473
rect 353298 151399 353354 151408
rect 229650 147656 229706 147665
rect 229650 147591 229652 147600
rect 229704 147591 229706 147600
rect 229652 147562 229704 147568
rect 3792 144900 3844 144906
rect 3792 144842 3844 144848
rect 230388 144900 230440 144906
rect 230388 144842 230440 144848
rect 353300 144900 353352 144906
rect 353300 144842 353352 144848
rect 230400 143857 230428 144842
rect 353312 144401 353340 144842
rect 353298 144392 353354 144401
rect 353298 144327 353354 144336
rect 230386 143848 230442 143857
rect 230386 143783 230442 143792
rect 353956 140865 353984 151778
rect 354048 147937 354076 178026
rect 354140 169289 354168 258062
rect 355336 209370 355364 456758
rect 356716 219366 356744 510614
rect 359476 230450 359504 563042
rect 360856 251190 360884 670686
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 367744 643136 367796 643142
rect 367744 643078 367796 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 364984 536852 365036 536858
rect 364984 536794 365036 536800
rect 363604 404388 363656 404394
rect 363604 404330 363656 404336
rect 360844 251184 360896 251190
rect 360844 251126 360896 251132
rect 359464 230444 359516 230450
rect 359464 230386 359516 230392
rect 356704 219360 356756 219366
rect 356704 219302 356756 219308
rect 355324 209364 355376 209370
rect 355324 209306 355376 209312
rect 363616 198694 363644 404330
rect 364996 226302 365024 536794
rect 367756 248402 367784 643078
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 374644 630692 374696 630698
rect 374644 630634 374696 630640
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 373264 524476 373316 524482
rect 373264 524418 373316 524424
rect 371884 430636 371936 430642
rect 371884 430578 371936 430584
rect 369124 324352 369176 324358
rect 369124 324294 369176 324300
rect 367744 248396 367796 248402
rect 367744 248338 367796 248344
rect 364984 226296 365036 226302
rect 364984 226238 365036 226244
rect 363604 198688 363656 198694
rect 363604 198630 363656 198636
rect 369136 183530 369164 324294
rect 371896 205630 371924 430578
rect 373276 223582 373304 524418
rect 374656 244254 374684 630634
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 381544 616888 381596 616894
rect 381544 616830 381596 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 378784 418192 378836 418198
rect 378784 418134 378836 418140
rect 377404 311908 377456 311914
rect 377404 311850 377456 311856
rect 374644 244248 374696 244254
rect 374644 244190 374696 244196
rect 373264 223576 373316 223582
rect 373264 223518 373316 223524
rect 371884 205624 371936 205630
rect 371884 205566 371936 205572
rect 369124 183524 369176 183530
rect 369124 183466 369176 183472
rect 377416 180810 377444 311850
rect 378796 201482 378824 418134
rect 381556 241466 381584 616830
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 580000 324358 580028 325207
rect 579988 324352 580040 324358
rect 579988 324294 580040 324300
rect 579802 312080 579858 312089
rect 579802 312015 579858 312024
rect 579816 311914 579844 312015
rect 579804 311908 579856 311914
rect 579804 311850 579856 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 442264 298172 442316 298178
rect 442264 298114 442316 298120
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 385684 244316 385736 244322
rect 385684 244258 385736 244264
rect 381544 241460 381596 241466
rect 381544 241402 381596 241408
rect 378784 201476 378836 201482
rect 378784 201418 378836 201424
rect 377404 180804 377456 180810
rect 377404 180746 377456 180752
rect 354126 169280 354182 169289
rect 354126 169215 354182 169224
rect 385696 167006 385724 244258
rect 442276 176662 442304 298114
rect 580276 259418 580304 697167
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580264 259412 580316 259418
rect 580264 259354 580316 259360
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 580368 237386 580396 590951
rect 580446 577688 580502 577697
rect 580446 577623 580502 577632
rect 580356 237380 580408 237386
rect 580356 237322 580408 237328
rect 580460 233238 580488 577623
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580448 233232 580500 233238
rect 580448 233174 580500 233180
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 442264 176656 442316 176662
rect 442264 176598 442316 176604
rect 385684 167000 385736 167006
rect 385684 166942 385736 166948
rect 580276 162858 580304 232319
rect 580552 219434 580580 484599
rect 580630 471472 580686 471481
rect 580630 471407 580686 471416
rect 580460 219406 580580 219434
rect 580460 216646 580488 219406
rect 580448 216640 580500 216646
rect 580448 216582 580500 216588
rect 580644 212498 580672 471407
rect 580722 378448 580778 378457
rect 580722 378383 580778 378392
rect 580632 212492 580684 212498
rect 580632 212434 580684 212440
rect 580354 205728 580410 205737
rect 580354 205663 580410 205672
rect 580264 162852 580316 162858
rect 580264 162794 580316 162800
rect 580368 155922 580396 205663
rect 580736 194546 580764 378383
rect 580814 351928 580870 351937
rect 580814 351863 580870 351872
rect 580724 194540 580776 194546
rect 580724 194482 580776 194488
rect 580446 192536 580502 192545
rect 580446 192471 580502 192480
rect 580356 155916 580408 155922
rect 580356 155858 580408 155864
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580184 151842 580212 152623
rect 580172 151836 580224 151842
rect 580172 151778 580224 151784
rect 580460 151774 580488 192471
rect 580828 187678 580856 351863
rect 580906 272232 580962 272241
rect 580906 272167 580962 272176
rect 580816 187672 580868 187678
rect 580816 187614 580868 187620
rect 580920 173874 580948 272167
rect 580908 173868 580960 173874
rect 580908 173810 580960 173816
rect 580538 165880 580594 165889
rect 580538 165815 580594 165824
rect 580448 151768 580500 151774
rect 580448 151710 580500 151716
rect 354034 147928 354090 147937
rect 354034 147863 354090 147872
rect 580552 144906 580580 165815
rect 580540 144900 580592 144906
rect 580540 144842 580592 144848
rect 353942 140856 353998 140865
rect 353942 140791 353998 140800
rect 3424 140752 3476 140758
rect 3424 140694 3476 140700
rect 230388 140752 230440 140758
rect 230388 140694 230440 140700
rect 230400 140049 230428 140694
rect 230386 140040 230442 140049
rect 230386 139975 230442 139984
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 353300 138032 353352 138038
rect 353300 137974 353352 137980
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 353312 137329 353340 137974
rect 353298 137320 353354 137329
rect 353298 137255 353354 137264
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3436 136610 3464 136711
rect 3424 136604 3476 136610
rect 3424 136546 3476 136552
rect 229836 136604 229888 136610
rect 229836 136546 229888 136552
rect 229848 136241 229876 136546
rect 229834 136232 229890 136241
rect 229834 136167 229890 136176
rect 354310 133784 354366 133793
rect 354310 133719 354366 133728
rect 229742 132424 229798 132433
rect 229742 132359 229798 132368
rect 3608 128376 3660 128382
rect 3608 128318 3660 128324
rect 3516 116000 3568 116006
rect 3516 115942 3568 115948
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3424 104916 3476 104922
rect 3424 104858 3476 104864
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 2780 49020 2832 49026
rect 2780 48962 2832 48968
rect 2792 6914 2820 48962
rect 3436 19417 3464 104858
rect 3528 58585 3556 115942
rect 3620 97617 3648 128318
rect 229756 111790 229784 132359
rect 353942 130248 353998 130257
rect 353942 130183 353998 130192
rect 230386 128616 230442 128625
rect 230386 128551 230442 128560
rect 230400 128382 230428 128551
rect 230388 128376 230440 128382
rect 230388 128318 230440 128324
rect 230110 124808 230166 124817
rect 230110 124743 230166 124752
rect 230018 121000 230074 121009
rect 230018 120935 230074 120944
rect 229926 113384 229982 113393
rect 229926 113319 229982 113328
rect 229744 111784 229796 111790
rect 229744 111726 229796 111732
rect 229834 109576 229890 109585
rect 229834 109511 229890 109520
rect 229742 101960 229798 101969
rect 229742 101895 229798 101904
rect 225604 97980 225656 97986
rect 225604 97922 225656 97928
rect 224316 97776 224368 97782
rect 224316 97718 224368 97724
rect 221464 97708 221516 97714
rect 221464 97650 221516 97656
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 124220 97436 124272 97442
rect 124220 97378 124272 97384
rect 106280 97368 106332 97374
rect 106280 97310 106332 97316
rect 10324 97300 10376 97306
rect 10324 97242 10376 97248
rect 4804 95940 4856 95946
rect 4804 95882 4856 95888
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2884 16574 2912 17206
rect 2884 16546 3648 16574
rect 2792 6886 2912 6914
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3324 1728 3330
rect 1676 3266 1728 3272
rect 1688 480 1716 3266
rect 2884 480 2912 6886
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 4816 3534 4844 95882
rect 7564 76560 7616 76566
rect 7564 76502 7616 76508
rect 6920 39364 6972 39370
rect 6920 39306 6972 39312
rect 6932 16574 6960 39306
rect 6932 16546 7512 16574
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 7484 3482 7512 16546
rect 7576 3602 7604 76502
rect 8300 51740 8352 51746
rect 8300 51682 8352 51688
rect 8312 16574 8340 51682
rect 8312 16546 8800 16574
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 5276 480 5304 3470
rect 7484 3454 7696 3482
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 9680 10328 9732 10334
rect 9680 10270 9732 10276
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 10270
rect 10336 3670 10364 97242
rect 80060 96008 80112 96014
rect 80060 95950 80112 95956
rect 60740 94512 60792 94518
rect 60740 94454 60792 94460
rect 46940 91792 46992 91798
rect 46940 91734 46992 91740
rect 26240 90364 26292 90370
rect 26240 90306 26292 90312
rect 16580 89004 16632 89010
rect 16580 88946 16632 88952
rect 13820 79348 13872 79354
rect 13820 79290 13872 79296
rect 11060 61396 11112 61402
rect 11060 61338 11112 61344
rect 11072 16574 11100 61338
rect 12440 60036 12492 60042
rect 12440 59978 12492 59984
rect 12452 16574 12480 59978
rect 13832 16574 13860 79290
rect 16592 16574 16620 88946
rect 20720 86284 20772 86290
rect 20720 86226 20772 86232
rect 17960 35216 18012 35222
rect 17960 35158 18012 35164
rect 11072 16546 11928 16574
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15948 480 15976 3470
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 35158
rect 20732 16574 20760 86226
rect 22100 36576 22152 36582
rect 22100 36518 22152 36524
rect 22112 16574 22140 36518
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19444 480 19472 3606
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20640 480 20668 3538
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24228 480 24256 3674
rect 25332 480 25360 3742
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 90306
rect 41420 76628 41472 76634
rect 41420 76570 41472 76576
rect 40040 75200 40092 75206
rect 40040 75142 40092 75148
rect 35900 73840 35952 73846
rect 35900 73782 35952 73788
rect 29000 72480 29052 72486
rect 29000 72422 29052 72428
rect 27620 24132 27672 24138
rect 27620 24074 27672 24080
rect 27632 16574 27660 24074
rect 29012 16574 29040 72422
rect 33140 46232 33192 46238
rect 33140 46174 33192 46180
rect 30380 19984 30432 19990
rect 30380 19926 30432 19932
rect 30392 16574 30420 19926
rect 33152 16574 33180 46174
rect 35912 16574 35940 73782
rect 40052 16574 40080 75142
rect 41432 16574 41460 76570
rect 44180 65544 44232 65550
rect 44180 65486 44232 65492
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 33152 16546 33640 16574
rect 35912 16546 36768 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 27724 480 27752 16546
rect 28908 3868 28960 3874
rect 28908 3810 28960 3816
rect 28920 480 28948 3810
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 32416 480 32444 3878
rect 33612 480 33640 16546
rect 34796 4820 34848 4826
rect 34796 4762 34848 4768
rect 34808 480 34836 4762
rect 35992 4004 36044 4010
rect 35992 3946 36044 3952
rect 36004 480 36032 3946
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 8968 38436 8974
rect 38384 8910 38436 8916
rect 38396 480 38424 8910
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 39592 480 39620 4014
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 43088 480 43116 4082
rect 44192 3398 44220 65486
rect 44272 40724 44324 40730
rect 44272 40666 44324 40672
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44284 480 44312 40666
rect 46952 16574 46980 91734
rect 53840 79416 53892 79422
rect 53840 79358 53892 79364
rect 48320 43444 48372 43450
rect 48320 43386 48372 43392
rect 48332 16574 48360 43386
rect 52460 42084 52512 42090
rect 52460 42026 52512 42032
rect 49700 18624 49752 18630
rect 49700 18566 49752 18572
rect 49712 16574 49740 18566
rect 52472 16574 52500 42026
rect 53852 16574 53880 79358
rect 57980 64184 58032 64190
rect 57980 64126 58032 64132
rect 56600 28280 56652 28286
rect 56600 28222 56652 28228
rect 55220 26920 55272 26926
rect 55220 26862 55272 26868
rect 55232 16574 55260 26862
rect 56612 16574 56640 28222
rect 57992 16574 58020 64126
rect 59360 47592 59412 47598
rect 59360 47534 59412 47540
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 52472 16546 52592 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 3334
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 7608 51408 7614
rect 51356 7550 51408 7556
rect 51368 480 51396 7550
rect 52564 480 52592 16546
rect 53288 14476 53340 14482
rect 53288 14418 53340 14424
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 14418
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 47534
rect 60752 3330 60780 94454
rect 71780 93152 71832 93158
rect 71780 93094 71832 93100
rect 69020 66904 69072 66910
rect 69020 66846 69072 66852
rect 64880 62824 64932 62830
rect 64880 62766 64932 62772
rect 63500 61464 63552 61470
rect 63500 61406 63552 61412
rect 62120 55888 62172 55894
rect 62120 55830 62172 55836
rect 60832 44872 60884 44878
rect 60832 44814 60884 44820
rect 60740 3324 60792 3330
rect 60740 3266 60792 3272
rect 60844 480 60872 44814
rect 62132 16574 62160 55830
rect 63512 16574 63540 61406
rect 64892 16574 64920 62766
rect 66260 50380 66312 50386
rect 66260 50322 66312 50328
rect 66272 16574 66300 50322
rect 67640 39432 67692 39438
rect 67640 39374 67692 39380
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3324 61712 3330
rect 61660 3266 61712 3272
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3266
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 39374
rect 69032 16574 69060 66846
rect 71792 16574 71820 93094
rect 78680 80708 78732 80714
rect 78680 80650 78732 80656
rect 74540 62892 74592 62898
rect 74540 62834 74592 62840
rect 73160 57248 73212 57254
rect 73160 57190 73212 57196
rect 73172 16574 73200 57190
rect 74552 16574 74580 62834
rect 77300 54528 77352 54534
rect 77300 54470 77352 54476
rect 77312 16574 77340 54470
rect 78692 16574 78720 80650
rect 80072 16574 80100 95950
rect 103520 87644 103572 87650
rect 103520 87586 103572 87592
rect 85580 83496 85632 83502
rect 85580 83438 85632 83444
rect 82820 65612 82872 65618
rect 82820 65554 82872 65560
rect 81440 40792 81492 40798
rect 81440 40734 81492 40740
rect 81452 16574 81480 40734
rect 82832 16574 82860 65554
rect 84200 58676 84252 58682
rect 84200 58618 84252 58624
rect 69032 16546 69152 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 77312 16546 77432 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 69124 480 69152 16546
rect 69848 15904 69900 15910
rect 69848 15846 69900 15852
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 15846
rect 71504 11756 71556 11762
rect 71504 11698 71556 11704
rect 71516 480 71544 11698
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 75920 11824 75972 11830
rect 75920 11766 75972 11772
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 11766
rect 77404 480 77432 16546
rect 78588 6180 78640 6186
rect 78588 6122 78640 6128
rect 78600 480 78628 6122
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 58618
rect 85592 3330 85620 83438
rect 89720 82136 89772 82142
rect 89720 82078 89772 82084
rect 88340 64252 88392 64258
rect 88340 64194 88392 64200
rect 86960 25560 87012 25566
rect 86960 25502 87012 25508
rect 85672 17332 85724 17338
rect 85672 17274 85724 17280
rect 85580 3324 85632 3330
rect 85580 3266 85632 3272
rect 85684 480 85712 17274
rect 86972 16574 87000 25502
rect 88352 16574 88380 64194
rect 89732 16574 89760 82078
rect 100760 77988 100812 77994
rect 100760 77930 100812 77936
rect 93860 68332 93912 68338
rect 93860 68274 93912 68280
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 86500 3324 86552 3330
rect 86500 3266 86552 3272
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3266
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 13116 91612 13122
rect 91560 13058 91612 13064
rect 91572 480 91600 13058
rect 92756 7676 92808 7682
rect 92756 7618 92808 7624
rect 92768 480 92796 7618
rect 93872 6914 93900 68274
rect 95240 66972 95292 66978
rect 95240 66914 95292 66920
rect 93952 22772 94004 22778
rect 93952 22714 94004 22720
rect 93964 16574 93992 22714
rect 95252 16574 95280 66914
rect 99380 46300 99432 46306
rect 99380 46242 99432 46248
rect 98000 33788 98052 33794
rect 98000 33730 98052 33736
rect 96620 28348 96672 28354
rect 96620 28290 96672 28296
rect 96632 16574 96660 28290
rect 98012 16574 98040 33730
rect 99392 16574 99420 46242
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 77930
rect 102140 37936 102192 37942
rect 102140 37878 102192 37884
rect 102152 6914 102180 37878
rect 102232 26988 102284 26994
rect 102232 26930 102284 26936
rect 102244 16574 102272 26930
rect 103532 16574 103560 87586
rect 104900 29640 104952 29646
rect 104900 29582 104952 29588
rect 104912 16574 104940 29582
rect 106292 16574 106320 97310
rect 113180 91860 113232 91866
rect 113180 91802 113232 91808
rect 107660 84856 107712 84862
rect 107660 84798 107712 84804
rect 107672 16574 107700 84798
rect 110420 69692 110472 69698
rect 110420 69634 110472 69640
rect 109040 31068 109092 31074
rect 109040 31010 109092 31016
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 31010
rect 110432 3330 110460 69634
rect 111800 49088 111852 49094
rect 111800 49030 111852 49036
rect 110512 42152 110564 42158
rect 110512 42094 110564 42100
rect 110420 3324 110472 3330
rect 110420 3266 110472 3272
rect 110524 480 110552 42094
rect 111812 16574 111840 49030
rect 113192 16574 113220 91802
rect 121460 71052 121512 71058
rect 121460 70994 121512 71000
rect 114560 53100 114612 53106
rect 114560 53042 114612 53048
rect 114572 16574 114600 53042
rect 118700 32428 118752 32434
rect 118700 32370 118752 32376
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 111616 3324 111668 3330
rect 111616 3266 111668 3272
rect 111628 480 111656 3266
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116400 14544 116452 14550
rect 116400 14486 116452 14492
rect 116412 480 116440 14486
rect 118712 3330 118740 32370
rect 118792 18692 118844 18698
rect 118792 18634 118844 18640
rect 118700 3324 118752 3330
rect 118700 3266 118752 3272
rect 117596 3256 117648 3262
rect 117596 3198 117648 3204
rect 117608 480 117636 3198
rect 118804 480 118832 18634
rect 121472 16574 121500 70994
rect 122840 21412 122892 21418
rect 122840 21354 122892 21360
rect 122852 16574 122880 21354
rect 124232 16574 124260 97378
rect 209780 96212 209832 96218
rect 209780 96154 209832 96160
rect 201500 96144 201552 96150
rect 201500 96086 201552 96092
rect 182180 96076 182232 96082
rect 182180 96018 182232 96024
rect 125600 94580 125652 94586
rect 125600 94522 125652 94528
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 119896 3324 119948 3330
rect 119896 3266 119948 3272
rect 119908 480 119936 3266
rect 121092 3256 121144 3262
rect 121092 3198 121144 3204
rect 121104 480 121132 3198
rect 122300 480 122328 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 94522
rect 160100 93220 160152 93226
rect 160100 93162 160152 93168
rect 151820 90432 151872 90438
rect 151820 90374 151872 90380
rect 147680 89072 147732 89078
rect 147680 89014 147732 89020
rect 139400 87712 139452 87718
rect 139400 87654 139452 87660
rect 126980 83564 127032 83570
rect 126980 83506 127032 83512
rect 126992 480 127020 83506
rect 129740 82204 129792 82210
rect 129740 82146 129792 82152
rect 128360 80776 128412 80782
rect 128360 80718 128412 80724
rect 127072 54596 127124 54602
rect 127072 54538 127124 54544
rect 127084 16574 127112 54538
rect 128372 16574 128400 80718
rect 129752 16574 129780 82146
rect 132500 78056 132552 78062
rect 132500 77998 132552 78004
rect 131120 58744 131172 58750
rect 131120 58686 131172 58692
rect 131132 16574 131160 58686
rect 132512 16574 132540 77998
rect 135260 75268 135312 75274
rect 135260 75210 135312 75216
rect 133880 57316 133932 57322
rect 133880 57258 133932 57264
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 57258
rect 135272 4214 135300 75210
rect 135352 38004 135404 38010
rect 135352 37946 135404 37952
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 135364 3482 135392 37946
rect 138020 36644 138072 36650
rect 138020 36586 138072 36592
rect 138032 16574 138060 36586
rect 139412 16574 139440 87654
rect 146300 86352 146352 86358
rect 146300 86294 146352 86300
rect 143540 73908 143592 73914
rect 143540 73850 143592 73856
rect 142160 35284 142212 35290
rect 142160 35226 142212 35232
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 137652 9036 137704 9042
rect 137652 8978 137704 8984
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 4150
rect 137664 480 137692 8978
rect 138860 480 138888 16546
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141240 10396 141292 10402
rect 141240 10338 141292 10344
rect 141252 480 141280 10338
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 35226
rect 143552 480 143580 73850
rect 143632 55956 143684 55962
rect 143632 55898 143684 55904
rect 143644 16574 143672 55898
rect 144920 20052 144972 20058
rect 144920 19994 144972 20000
rect 144932 16574 144960 19994
rect 146312 16574 146340 86294
rect 147692 16574 147720 89014
rect 150440 79484 150492 79490
rect 150440 79426 150492 79432
rect 149060 60104 149112 60110
rect 149060 60046 149112 60052
rect 149072 16574 149100 60046
rect 150452 16574 150480 79426
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 90374
rect 153200 72548 153252 72554
rect 153200 72490 153252 72496
rect 151912 33856 151964 33862
rect 151912 33798 151964 33804
rect 151924 16574 151952 33798
rect 153212 16574 153240 72490
rect 157340 69760 157392 69766
rect 157340 69702 157392 69708
rect 155960 31136 156012 31142
rect 155960 31078 156012 31084
rect 154580 24200 154632 24206
rect 154580 24142 154632 24148
rect 154592 16574 154620 24142
rect 155972 16574 156000 31078
rect 157352 16574 157380 69702
rect 158720 21480 158772 21486
rect 158720 21422 158772 21428
rect 158732 16574 158760 21422
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11694 160140 93162
rect 164240 91928 164292 91934
rect 164240 91870 164292 91876
rect 161480 68400 161532 68406
rect 161480 68342 161532 68348
rect 160192 29708 160244 29714
rect 160192 29650 160244 29656
rect 160100 11688 160152 11694
rect 160100 11630 160152 11636
rect 160204 6914 160232 29650
rect 161492 16574 161520 68342
rect 162860 53168 162912 53174
rect 162860 53110 162912 53116
rect 162872 16574 162900 53110
rect 164252 16574 164280 91870
rect 171140 90500 171192 90506
rect 171140 90442 171192 90448
rect 168380 76696 168432 76702
rect 168380 76638 168432 76644
rect 165620 67040 165672 67046
rect 165620 66982 165672 66988
rect 165632 16574 165660 66982
rect 167000 51808 167052 51814
rect 167000 51750 167052 51756
rect 167012 16574 167040 51750
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11688 161348 11694
rect 161296 11630 161348 11636
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11630
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 3194 168420 76638
rect 169760 50448 169812 50454
rect 169760 50390 169812 50396
rect 169772 16574 169800 50390
rect 171152 16574 171180 90442
rect 175280 89140 175332 89146
rect 175280 89082 175332 89088
rect 173900 75336 173952 75342
rect 173900 75278 173952 75284
rect 172520 65680 172572 65686
rect 172520 65622 172572 65628
rect 172532 16574 172560 65622
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 168472 4888 168524 4894
rect 168472 4830 168524 4836
rect 168380 3188 168432 3194
rect 168380 3130 168432 3136
rect 168484 2530 168512 4830
rect 169576 3188 169628 3194
rect 169576 3130 169628 3136
rect 168392 2502 168512 2530
rect 168392 480 168420 2502
rect 169588 480 169616 3130
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 75278
rect 175292 16574 175320 89082
rect 178040 87780 178092 87786
rect 178040 87722 178092 87728
rect 176660 47660 176712 47666
rect 176660 47602 176712 47608
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 11694 176700 47602
rect 176752 22840 176804 22846
rect 176752 22782 176804 22788
rect 176660 11688 176712 11694
rect 176660 11630 176712 11636
rect 176764 6914 176792 22782
rect 178052 16574 178080 87722
rect 180800 73976 180852 73982
rect 180800 73918 180852 73924
rect 179420 64320 179472 64326
rect 179420 64262 179472 64268
rect 179432 16574 179460 64262
rect 180812 16574 180840 73918
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 11688 177908 11694
rect 177856 11630 177908 11636
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177868 480 177896 11630
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 96018
rect 195980 94648 196032 94654
rect 195980 94590 196032 94596
rect 193220 93288 193272 93294
rect 193220 93230 193272 93236
rect 184940 86420 184992 86426
rect 184940 86362 184992 86368
rect 183560 62960 183612 62966
rect 183560 62902 183612 62908
rect 183572 16574 183600 62902
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11694 184980 86362
rect 189080 83632 189132 83638
rect 189080 83574 189132 83580
rect 186320 61532 186372 61538
rect 186320 61474 186372 61480
rect 185032 25628 185084 25634
rect 185032 25570 185084 25576
rect 184940 11688 184992 11694
rect 184940 11630 184992 11636
rect 185044 6914 185072 25570
rect 186332 16574 186360 61474
rect 187700 46368 187752 46374
rect 187700 46310 187752 46316
rect 187712 16574 187740 46310
rect 189092 16574 189120 83574
rect 191840 43512 191892 43518
rect 191840 43454 191892 43460
rect 191852 16574 191880 43454
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 191852 16546 192064 16574
rect 186136 11688 186188 11694
rect 186136 11630 186188 11636
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11630
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 190460 13184 190512 13190
rect 190460 13126 190512 13132
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 13126
rect 192036 480 192064 16546
rect 193232 4214 193260 93230
rect 193312 82272 193364 82278
rect 193312 82214 193364 82220
rect 193220 4208 193272 4214
rect 193220 4150 193272 4156
rect 193324 3482 193352 82214
rect 194600 42220 194652 42226
rect 194600 42162 194652 42168
rect 194612 16574 194640 42162
rect 195992 16574 196020 94590
rect 200120 93356 200172 93362
rect 200120 93298 200172 93304
rect 197360 78124 197412 78130
rect 197360 78066 197412 78072
rect 197372 16574 197400 78066
rect 198740 72616 198792 72622
rect 198740 72558 198792 72564
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194416 4208 194468 4214
rect 194416 4150 194468 4156
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 4150
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 72558
rect 200132 16574 200160 93298
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 11694 201540 96086
rect 207020 91996 207072 92002
rect 207020 91938 207072 91944
rect 202880 84924 202932 84930
rect 202880 84866 202932 84872
rect 201592 71120 201644 71126
rect 201592 71062 201644 71068
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 71062
rect 202892 16574 202920 84866
rect 205640 40860 205692 40866
rect 205640 40802 205692 40808
rect 205652 16574 205680 40802
rect 202892 16546 203472 16574
rect 205652 16546 206232 16574
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205088 15972 205140 15978
rect 205088 15914 205140 15920
rect 205100 480 205128 15914
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 91938
rect 208400 60172 208452 60178
rect 208400 60114 208452 60120
rect 208412 16574 208440 60114
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 96154
rect 215300 92064 215352 92070
rect 215300 92006 215352 92012
rect 213920 90568 213972 90574
rect 213920 90510 213972 90516
rect 211160 80844 211212 80850
rect 211160 80786 211212 80792
rect 209872 69828 209924 69834
rect 209872 69770 209924 69776
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 69770
rect 211172 16574 211200 80786
rect 212540 27056 212592 27062
rect 212540 26998 212592 27004
rect 212552 16574 212580 26998
rect 213932 16574 213960 90510
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 92006
rect 220820 89208 220872 89214
rect 220820 89150 220872 89156
rect 219440 86488 219492 86494
rect 219440 86430 219492 86436
rect 218060 84992 218112 84998
rect 218060 84934 218112 84940
rect 216680 68468 216732 68474
rect 216680 68410 216732 68416
rect 216692 16574 216720 68410
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 4214 218100 84934
rect 219452 16574 219480 86430
rect 220832 16574 220860 89150
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 218152 7744 218204 7750
rect 218152 7686 218204 7692
rect 218060 4208 218112 4214
rect 218060 4150 218112 4156
rect 218164 3482 218192 7686
rect 219256 4208 219308 4214
rect 219256 4150 219308 4156
rect 218072 3454 218192 3482
rect 218072 480 218100 3454
rect 219268 480 219296 4150
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 221476 7614 221504 97650
rect 224224 97640 224276 97646
rect 224224 97582 224276 97588
rect 222200 58812 222252 58818
rect 222200 58754 222252 58760
rect 222212 16574 222240 58754
rect 223580 39500 223632 39506
rect 223580 39442 223632 39448
rect 222212 16546 222792 16574
rect 221464 7608 221516 7614
rect 221464 7550 221516 7556
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 39442
rect 224236 9042 224264 97582
rect 224328 40730 224356 97718
rect 224960 79552 225012 79558
rect 224960 79494 225012 79500
rect 224316 40724 224368 40730
rect 224316 40666 224368 40672
rect 224972 16574 225000 79494
rect 224972 16546 225184 16574
rect 224224 9036 224276 9042
rect 224224 8978 224276 8984
rect 225156 480 225184 16546
rect 225616 7750 225644 97922
rect 228364 97572 228416 97578
rect 228364 97514 228416 97520
rect 227720 94716 227772 94722
rect 227720 94658 227772 94664
rect 226340 44940 226392 44946
rect 226340 44882 226392 44888
rect 226352 11694 226380 44882
rect 226432 17400 226484 17406
rect 226432 17342 226484 17348
rect 226340 11688 226392 11694
rect 226340 11630 226392 11636
rect 225604 7744 225656 7750
rect 225604 7686 225656 7692
rect 226444 6914 226472 17342
rect 227732 16574 227760 94658
rect 227732 16546 228312 16574
rect 227536 11688 227588 11694
rect 227536 11630 227588 11636
rect 226352 6886 226472 6914
rect 226352 480 226380 6886
rect 227548 480 227576 11630
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228376 4894 228404 97514
rect 229100 49156 229152 49162
rect 229100 49098 229152 49104
rect 229112 16574 229140 49098
rect 229112 16546 229416 16574
rect 228364 4888 228416 4894
rect 228364 4830 228416 4836
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 229756 6866 229784 101895
rect 229848 33114 229876 109511
rect 229940 45558 229968 113319
rect 230032 71738 230060 120935
rect 230124 85542 230152 124743
rect 230202 117192 230258 117201
rect 230202 117127 230258 117136
rect 230216 116006 230244 117127
rect 230204 116000 230256 116006
rect 230204 115942 230256 115948
rect 353956 113150 353984 130183
rect 354324 126954 354352 133719
rect 354312 126948 354364 126954
rect 354312 126890 354364 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 354586 126576 354642 126585
rect 354586 126511 354642 126520
rect 354494 123040 354550 123049
rect 354494 122975 354550 122984
rect 354402 119504 354458 119513
rect 354402 119439 354458 119448
rect 354310 115968 354366 115977
rect 354310 115903 354366 115912
rect 353944 113144 353996 113150
rect 353944 113086 353996 113092
rect 354218 112432 354274 112441
rect 354218 112367 354274 112376
rect 354126 108896 354182 108905
rect 354126 108831 354182 108840
rect 230386 105768 230442 105777
rect 230386 105703 230442 105712
rect 230400 104922 230428 105703
rect 354034 105360 354090 105369
rect 354034 105295 354090 105304
rect 230388 104916 230440 104922
rect 230388 104858 230440 104864
rect 353942 101824 353998 101833
rect 353942 101759 353998 101768
rect 239232 100162 239430 100178
rect 285968 100162 286166 100178
rect 238760 100156 238812 100162
rect 238760 100098 238812 100104
rect 239220 100156 239430 100162
rect 239272 100150 239430 100156
rect 285680 100156 285732 100162
rect 239220 100098 239272 100104
rect 285680 100098 285732 100104
rect 285956 100156 286166 100162
rect 286008 100150 286166 100156
rect 285956 100098 286008 100104
rect 231124 97028 231176 97034
rect 231124 96970 231176 96976
rect 230480 87848 230532 87854
rect 230480 87790 230532 87796
rect 230112 85536 230164 85542
rect 230112 85478 230164 85484
rect 230020 71732 230072 71738
rect 230020 71674 230072 71680
rect 229928 45552 229980 45558
rect 229928 45494 229980 45500
rect 229836 33108 229888 33114
rect 229836 33050 229888 33056
rect 230492 16574 230520 87790
rect 231136 39370 231164 96970
rect 231952 96960 232004 96966
rect 231952 96902 232004 96908
rect 231860 76764 231912 76770
rect 231860 76706 231912 76712
rect 231124 39364 231176 39370
rect 231124 39306 231176 39312
rect 230492 16546 231072 16574
rect 229744 6860 229796 6866
rect 229744 6802 229796 6808
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 76706
rect 231964 17270 231992 96902
rect 232148 95946 232176 100028
rect 232136 95940 232188 95946
rect 232136 95882 232188 95888
rect 232332 84194 232360 100028
rect 232504 96756 232556 96762
rect 232504 96698 232556 96704
rect 232240 84166 232360 84194
rect 232240 76566 232268 84166
rect 232228 76560 232280 76566
rect 232228 76502 232280 76508
rect 232516 61402 232544 96698
rect 232504 61396 232556 61402
rect 232504 61338 232556 61344
rect 232608 49026 232636 100028
rect 232792 96966 232820 100028
rect 233068 97306 233096 100028
rect 233056 97300 233108 97306
rect 233056 97242 233108 97248
rect 232780 96960 232832 96966
rect 232780 96902 232832 96908
rect 232596 49020 232648 49026
rect 232596 48962 232648 48968
rect 231952 17264 232004 17270
rect 231952 17206 232004 17212
rect 233344 3369 233372 100028
rect 233528 97034 233556 100028
rect 233516 97028 233568 97034
rect 233516 96970 233568 96976
rect 233608 96960 233660 96966
rect 233608 96902 233660 96908
rect 233424 7608 233476 7614
rect 233424 7550 233476 7556
rect 233330 3360 233386 3369
rect 233330 3295 233386 3304
rect 233436 480 233464 7550
rect 233620 3466 233648 96902
rect 233804 84194 233832 100028
rect 233884 97028 233936 97034
rect 233884 96970 233936 96976
rect 233896 86290 233924 96970
rect 233884 86284 233936 86290
rect 233884 86226 233936 86232
rect 234080 84194 234108 100028
rect 234264 96966 234292 100028
rect 234252 96960 234304 96966
rect 234252 96902 234304 96908
rect 234540 96762 234568 100028
rect 234620 96960 234672 96966
rect 234620 96902 234672 96908
rect 234528 96756 234580 96762
rect 234528 96698 234580 96704
rect 234632 89010 234660 96902
rect 234620 89004 234672 89010
rect 234620 88946 234672 88952
rect 233712 84166 233832 84194
rect 233988 84166 234108 84194
rect 233712 51746 233740 84166
rect 233700 51740 233752 51746
rect 233700 51682 233752 51688
rect 233988 10334 234016 84166
rect 234816 60042 234844 100028
rect 235000 84194 235028 100028
rect 234908 84166 235028 84194
rect 235092 100014 235290 100042
rect 235368 100014 235566 100042
rect 234908 79354 234936 84166
rect 234896 79348 234948 79354
rect 234896 79290 234948 79296
rect 234804 60036 234856 60042
rect 234804 59978 234856 59984
rect 233976 10328 234028 10334
rect 233976 10270 234028 10276
rect 234620 10328 234672 10334
rect 234620 10270 234672 10276
rect 233608 3460 233660 3466
rect 233608 3402 233660 3408
rect 234632 480 234660 10270
rect 235092 3534 235120 100014
rect 235368 96966 235396 100014
rect 235356 96960 235408 96966
rect 235356 96902 235408 96908
rect 235264 96892 235316 96898
rect 235264 96834 235316 96840
rect 235276 36582 235304 96834
rect 235736 84194 235764 100028
rect 235368 84166 235764 84194
rect 235264 36576 235316 36582
rect 235264 36518 235316 36524
rect 235368 35222 235396 84166
rect 235356 35216 235408 35222
rect 235356 35158 235408 35164
rect 235816 4888 235868 4894
rect 235816 4830 235868 4836
rect 235080 3528 235132 3534
rect 235080 3470 235132 3476
rect 235828 480 235856 4830
rect 236012 3670 236040 100028
rect 236210 100014 236316 100042
rect 236000 3664 236052 3670
rect 236000 3606 236052 3612
rect 236288 3602 236316 100014
rect 236472 97034 236500 100028
rect 236460 97028 236512 97034
rect 236460 96970 236512 96976
rect 236748 96898 236776 100028
rect 236736 96892 236788 96898
rect 236736 96834 236788 96840
rect 236932 84194 236960 100028
rect 236840 84166 236960 84194
rect 237024 100014 237222 100042
rect 236840 3738 236868 84166
rect 237024 6914 237052 100014
rect 237484 90370 237512 100028
rect 237472 90364 237524 90370
rect 237472 90306 237524 90312
rect 237668 24138 237696 100028
rect 237748 96960 237800 96966
rect 237748 96902 237800 96908
rect 237760 72486 237788 96902
rect 237944 84194 237972 100028
rect 238036 100014 238234 100042
rect 238036 96966 238064 100014
rect 238024 96960 238076 96966
rect 238024 96902 238076 96908
rect 238024 96824 238076 96830
rect 238024 96766 238076 96772
rect 237852 84166 237972 84194
rect 237748 72480 237800 72486
rect 237748 72422 237800 72428
rect 237656 24132 237708 24138
rect 237656 24074 237708 24080
rect 236932 6886 237052 6914
rect 236932 3806 236960 6886
rect 237012 4956 237064 4962
rect 237012 4898 237064 4904
rect 236920 3800 236972 3806
rect 236920 3742 236972 3748
rect 236828 3732 236880 3738
rect 236828 3674 236880 3680
rect 236276 3596 236328 3602
rect 236276 3538 236328 3544
rect 237024 480 237052 4898
rect 237852 3874 237880 84166
rect 238036 3942 238064 96766
rect 238404 84194 238432 100028
rect 238496 100014 238694 100042
rect 238496 96830 238524 100014
rect 238484 96824 238536 96830
rect 238484 96766 238536 96772
rect 238312 84166 238432 84194
rect 238312 19990 238340 84166
rect 238300 19984 238352 19990
rect 238300 19926 238352 19932
rect 238116 9036 238168 9042
rect 238116 8978 238168 8984
rect 238024 3936 238076 3942
rect 238024 3878 238076 3884
rect 237840 3868 237892 3874
rect 237840 3810 237892 3816
rect 238128 480 238156 8978
rect 238772 4010 238800 100098
rect 238956 84194 238984 100028
rect 239154 100014 239260 100042
rect 238864 84166 238984 84194
rect 238864 46238 238892 84166
rect 238852 46232 238904 46238
rect 238852 46174 238904 46180
rect 239232 4826 239260 100014
rect 239404 96960 239456 96966
rect 239404 96902 239456 96908
rect 239416 75206 239444 96902
rect 239600 84194 239628 100028
rect 239508 84166 239628 84194
rect 239692 100014 239890 100042
rect 239404 75200 239456 75206
rect 239404 75142 239456 75148
rect 239508 73846 239536 84166
rect 239496 73840 239548 73846
rect 239496 73782 239548 73788
rect 239692 8974 239720 100014
rect 240152 96898 240180 100028
rect 240336 96966 240364 100028
rect 240428 100014 240626 100042
rect 240704 100014 240902 100042
rect 240324 96960 240376 96966
rect 240324 96902 240376 96908
rect 240140 96892 240192 96898
rect 240140 96834 240192 96840
rect 240428 76634 240456 100014
rect 240416 76628 240468 76634
rect 240416 76570 240468 76576
rect 239680 8968 239732 8974
rect 239680 8910 239732 8916
rect 239312 6384 239364 6390
rect 239312 6326 239364 6332
rect 239220 4820 239272 4826
rect 239220 4762 239272 4768
rect 238760 4004 238812 4010
rect 238760 3946 238812 3952
rect 239324 480 239352 6326
rect 240508 6248 240560 6254
rect 240508 6190 240560 6196
rect 240520 480 240548 6190
rect 240704 4146 240732 100014
rect 241072 97782 241100 100028
rect 241060 97776 241112 97782
rect 241060 97718 241112 97724
rect 241348 84194 241376 100028
rect 241428 96892 241480 96898
rect 241428 96834 241480 96840
rect 241256 84166 241376 84194
rect 241256 65550 241284 84166
rect 241244 65544 241296 65550
rect 241244 65486 241296 65492
rect 240692 4140 240744 4146
rect 240692 4082 240744 4088
rect 241440 4078 241468 96834
rect 241624 84194 241652 100028
rect 241822 100014 241928 100042
rect 241900 91798 241928 100014
rect 241888 91792 241940 91798
rect 241888 91734 241940 91740
rect 242084 84194 242112 100028
rect 242164 96960 242216 96966
rect 242164 96902 242216 96908
rect 241532 84166 241652 84194
rect 241992 84166 242112 84194
rect 241428 4072 241480 4078
rect 241428 4014 241480 4020
rect 241532 3398 241560 84166
rect 241992 43450 242020 84166
rect 242176 62830 242204 96902
rect 242360 84194 242388 100028
rect 242544 97714 242572 100028
rect 242636 100014 242834 100042
rect 242912 100014 243110 100042
rect 242532 97708 242584 97714
rect 242532 97650 242584 97656
rect 242268 84166 242388 84194
rect 242164 62824 242216 62830
rect 242164 62766 242216 62772
rect 241980 43444 242032 43450
rect 241980 43386 242032 43392
rect 242268 18630 242296 84166
rect 242636 42090 242664 100014
rect 242624 42084 242676 42090
rect 242624 42026 242676 42032
rect 242256 18624 242308 18630
rect 242256 18566 242308 18572
rect 242912 14482 242940 100014
rect 242992 97096 243044 97102
rect 242992 97038 243044 97044
rect 243004 94518 243032 97038
rect 242992 94512 243044 94518
rect 242992 94454 243044 94460
rect 243280 79422 243308 100028
rect 243556 96914 243584 100028
rect 243360 96892 243412 96898
rect 243360 96834 243412 96840
rect 243464 96886 243584 96914
rect 243740 96898 243768 100028
rect 243832 100014 244030 100042
rect 243728 96892 243780 96898
rect 243268 79416 243320 79422
rect 243268 79358 243320 79364
rect 243372 28286 243400 96834
rect 243360 28280 243412 28286
rect 243360 28222 243412 28228
rect 243464 26926 243492 96886
rect 243728 96834 243780 96840
rect 243544 96824 243596 96830
rect 243544 96766 243596 96772
rect 243556 47598 243584 96766
rect 243832 64190 243860 100014
rect 244292 96830 244320 100028
rect 244490 100014 244596 100042
rect 244280 96824 244332 96830
rect 244280 96766 244332 96772
rect 243820 64184 243872 64190
rect 243820 64126 243872 64132
rect 243544 47592 243596 47598
rect 243544 47534 243596 47540
rect 244568 44878 244596 100014
rect 244752 97102 244780 100028
rect 244844 100014 245042 100042
rect 244740 97096 244792 97102
rect 244740 97038 244792 97044
rect 244844 55894 244872 100014
rect 245212 84194 245240 100028
rect 245488 96966 245516 100028
rect 245476 96960 245528 96966
rect 245476 96902 245528 96908
rect 245120 84166 245240 84194
rect 245120 61470 245148 84166
rect 245108 61464 245160 61470
rect 245108 61406 245160 61412
rect 244832 55888 244884 55894
rect 244832 55830 244884 55836
rect 245764 50386 245792 100028
rect 245948 84194 245976 100028
rect 245856 84166 245976 84194
rect 246040 100014 246238 100042
rect 245752 50380 245804 50386
rect 245752 50322 245804 50328
rect 244556 44872 244608 44878
rect 244556 44814 244608 44820
rect 245856 39438 245884 84166
rect 246040 66910 246068 100014
rect 246304 94512 246356 94518
rect 246304 94454 246356 94460
rect 246028 66904 246080 66910
rect 246028 66846 246080 66852
rect 245844 39432 245896 39438
rect 245844 39374 245896 39380
rect 243452 26920 243504 26926
rect 243452 26862 243504 26868
rect 242992 18624 243044 18630
rect 242992 18566 243044 18572
rect 243004 16574 243032 18566
rect 243004 16546 244136 16574
rect 242900 14476 242952 14482
rect 242900 14418 242952 14424
rect 241704 7812 241756 7818
rect 241704 7754 241756 7760
rect 241520 3392 241572 3398
rect 241520 3334 241572 3340
rect 241716 480 241744 7754
rect 242900 7744 242952 7750
rect 242900 7686 242952 7692
rect 242912 480 242940 7686
rect 244108 480 244136 16546
rect 246316 11762 246344 94454
rect 246500 89714 246528 100028
rect 246684 94518 246712 100028
rect 246776 100014 246974 100042
rect 246672 94512 246724 94518
rect 246672 94454 246724 94460
rect 246776 93158 246804 100014
rect 246764 93152 246816 93158
rect 246764 93094 246816 93100
rect 246408 89686 246528 89714
rect 246408 15910 246436 89686
rect 247144 84194 247172 100028
rect 247224 94444 247276 94450
rect 247224 94386 247276 94392
rect 247052 84166 247172 84194
rect 247052 57254 247080 84166
rect 247040 57248 247092 57254
rect 247040 57190 247092 57196
rect 247236 54534 247264 94386
rect 247420 62898 247448 100028
rect 247696 99374 247724 100028
rect 247604 99346 247724 99374
rect 247500 94512 247552 94518
rect 247500 94454 247552 94460
rect 247408 62892 247460 62898
rect 247408 62834 247460 62840
rect 247224 54528 247276 54534
rect 247224 54470 247276 54476
rect 246396 15904 246448 15910
rect 246396 15846 246448 15852
rect 246304 11756 246356 11762
rect 246304 11698 246356 11704
rect 247408 11756 247460 11762
rect 247408 11698 247460 11704
rect 246396 8968 246448 8974
rect 246396 8910 246448 8916
rect 245200 4820 245252 4826
rect 245200 4762 245252 4768
rect 245212 480 245240 4762
rect 246408 480 246436 8910
rect 247420 3482 247448 11698
rect 247512 6186 247540 94454
rect 247604 11830 247632 99346
rect 247684 96688 247736 96694
rect 247684 96630 247736 96636
rect 247696 80714 247724 96630
rect 247880 94450 247908 100028
rect 247972 100014 248170 100042
rect 247972 94518 248000 100014
rect 248432 96694 248460 100028
rect 248420 96688 248472 96694
rect 248420 96630 248472 96636
rect 248616 96014 248644 100028
rect 248604 96008 248656 96014
rect 248604 95950 248656 95956
rect 247960 94512 248012 94518
rect 247960 94454 248012 94460
rect 248696 94512 248748 94518
rect 248696 94454 248748 94460
rect 247868 94444 247920 94450
rect 247868 94386 247920 94392
rect 247684 80708 247736 80714
rect 247684 80650 247736 80656
rect 248708 65618 248736 94454
rect 248892 84194 248920 100028
rect 248984 100014 249182 100042
rect 248984 94518 249012 100014
rect 248972 94512 249024 94518
rect 248972 94454 249024 94460
rect 248972 94376 249024 94382
rect 248972 94318 249024 94324
rect 248800 84166 248920 84194
rect 248696 65612 248748 65618
rect 248696 65554 248748 65560
rect 248800 40798 248828 84166
rect 248788 40792 248840 40798
rect 248788 40734 248840 40740
rect 248984 17338 249012 94318
rect 249352 84194 249380 100028
rect 249444 100014 249642 100042
rect 249444 94382 249472 100014
rect 249432 94376 249484 94382
rect 249432 94318 249484 94324
rect 249904 84194 249932 100028
rect 250088 84194 250116 100028
rect 250168 94512 250220 94518
rect 250168 94454 250220 94460
rect 249260 84166 249380 84194
rect 249812 84166 249932 84194
rect 249996 84166 250116 84194
rect 249260 58682 249288 84166
rect 249812 83502 249840 84166
rect 249800 83496 249852 83502
rect 249800 83438 249852 83444
rect 249248 58676 249300 58682
rect 249248 58618 249300 58624
rect 249996 25566 250024 84166
rect 250180 82142 250208 94454
rect 250364 84194 250392 100028
rect 250456 100014 250654 100042
rect 250456 94518 250484 100014
rect 250444 94512 250496 94518
rect 250444 94454 250496 94460
rect 250444 94376 250496 94382
rect 250444 94318 250496 94324
rect 250272 84166 250392 84194
rect 250168 82136 250220 82142
rect 250168 82078 250220 82084
rect 250272 64258 250300 84166
rect 250260 64252 250312 64258
rect 250260 64194 250312 64200
rect 249984 25560 250036 25566
rect 249984 25502 250036 25508
rect 248972 17332 249024 17338
rect 248972 17274 249024 17280
rect 247592 11824 247644 11830
rect 247592 11766 247644 11772
rect 250456 7682 250484 94318
rect 250824 84194 250852 100028
rect 250916 100014 251114 100042
rect 250916 94382 250944 100014
rect 250904 94376 250956 94382
rect 250904 94318 250956 94324
rect 251284 84194 251312 100028
rect 251574 100014 251680 100042
rect 251364 94512 251416 94518
rect 251364 94454 251416 94460
rect 250732 84166 250852 84194
rect 251192 84166 251312 84194
rect 250732 13122 250760 84166
rect 251192 68338 251220 84166
rect 251180 68332 251232 68338
rect 251180 68274 251232 68280
rect 251376 33794 251404 94454
rect 251364 33788 251416 33794
rect 251364 33730 251416 33736
rect 251652 22778 251680 100014
rect 251836 84194 251864 100028
rect 252020 84194 252048 100028
rect 252112 100014 252310 100042
rect 252112 94518 252140 100014
rect 252572 94518 252600 100028
rect 252100 94512 252152 94518
rect 252100 94454 252152 94460
rect 252560 94512 252612 94518
rect 252560 94454 252612 94460
rect 252756 89714 252784 100028
rect 252836 94512 252888 94518
rect 252836 94454 252888 94460
rect 251744 84166 251864 84194
rect 251928 84166 252048 84194
rect 252664 89686 252784 89714
rect 251744 66978 251772 84166
rect 251732 66972 251784 66978
rect 251732 66914 251784 66920
rect 251928 28354 251956 84166
rect 252664 77994 252692 89686
rect 252652 77988 252704 77994
rect 252652 77930 252704 77936
rect 252848 46306 252876 94454
rect 252836 46300 252888 46306
rect 252836 46242 252888 46248
rect 253032 37942 253060 100028
rect 253124 100014 253322 100042
rect 253020 37936 253072 37942
rect 253020 37878 253072 37884
rect 251916 28348 251968 28354
rect 251916 28290 251968 28296
rect 253124 26994 253152 100014
rect 253492 87650 253520 100028
rect 253584 100014 253782 100042
rect 253480 87644 253532 87650
rect 253480 87586 253532 87592
rect 253584 29646 253612 100014
rect 254044 97374 254072 100028
rect 254242 100014 254348 100042
rect 254032 97368 254084 97374
rect 254032 97310 254084 97316
rect 254320 84862 254348 100014
rect 254308 84856 254360 84862
rect 254308 84798 254360 84804
rect 254504 84194 254532 100028
rect 254688 84194 254716 100028
rect 254412 84166 254532 84194
rect 254596 84166 254716 84194
rect 254780 100014 254978 100042
rect 255056 100014 255254 100042
rect 254412 31074 254440 84166
rect 254596 42158 254624 84166
rect 254780 69698 254808 100014
rect 254768 69692 254820 69698
rect 254768 69634 254820 69640
rect 255056 49094 255084 100014
rect 255424 91866 255452 100028
rect 255504 96892 255556 96898
rect 255504 96834 255556 96840
rect 255412 91860 255464 91866
rect 255412 91802 255464 91808
rect 255044 49088 255096 49094
rect 255044 49030 255096 49036
rect 254584 42152 254636 42158
rect 254584 42094 254636 42100
rect 254400 31068 254452 31074
rect 254400 31010 254452 31016
rect 253572 29640 253624 29646
rect 253572 29582 253624 29588
rect 253112 26988 253164 26994
rect 253112 26930 253164 26936
rect 251640 22772 251692 22778
rect 251640 22714 251692 22720
rect 255516 18698 255544 96834
rect 255700 84194 255728 100028
rect 255976 97866 256004 100028
rect 255884 97838 256004 97866
rect 255780 96960 255832 96966
rect 255780 96902 255832 96908
rect 255608 84166 255728 84194
rect 255608 53106 255636 84166
rect 255596 53100 255648 53106
rect 255596 53042 255648 53048
rect 255504 18692 255556 18698
rect 255504 18634 255556 18640
rect 251180 14476 251232 14482
rect 251180 14418 251232 14424
rect 250720 13116 250772 13122
rect 250720 13058 250772 13064
rect 250444 7676 250496 7682
rect 250444 7618 250496 7624
rect 247500 6180 247552 6186
rect 247500 6122 247552 6128
rect 248788 6180 248840 6186
rect 248788 6122 248840 6128
rect 247420 3454 247632 3482
rect 247604 480 247632 3454
rect 248800 480 248828 6122
rect 249984 5024 250036 5030
rect 249984 4966 250036 4972
rect 249996 480 250024 4966
rect 251192 480 251220 14418
rect 252376 13116 252428 13122
rect 252376 13058 252428 13064
rect 252388 480 252416 13058
rect 254676 9104 254728 9110
rect 254676 9046 254728 9052
rect 253480 6316 253532 6322
rect 253480 6258 253532 6264
rect 253492 480 253520 6258
rect 254688 480 254716 9046
rect 255792 3330 255820 96902
rect 255884 14550 255912 97838
rect 255964 97776 256016 97782
rect 255964 97718 256016 97724
rect 255976 78062 256004 97718
rect 256160 96966 256188 100028
rect 256252 100014 256450 100042
rect 256148 96960 256200 96966
rect 256148 96902 256200 96908
rect 256252 96898 256280 100014
rect 256240 96892 256292 96898
rect 256240 96834 256292 96840
rect 256712 93854 256740 100028
rect 256910 100014 257016 100042
rect 256988 96966 257016 100014
rect 257172 98002 257200 100028
rect 257080 97974 257200 98002
rect 256976 96960 257028 96966
rect 256976 96902 257028 96908
rect 256712 93826 257016 93854
rect 256792 80708 256844 80714
rect 256792 80650 256844 80656
rect 255964 78056 256016 78062
rect 255964 77998 256016 78004
rect 255872 14544 255924 14550
rect 255872 14486 255924 14492
rect 255872 3460 255924 3466
rect 255872 3402 255924 3408
rect 255780 3324 255832 3330
rect 255780 3266 255832 3272
rect 255884 480 255912 3402
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256804 354 256832 80650
rect 256988 32434 257016 93826
rect 257080 71058 257108 97974
rect 257160 97912 257212 97918
rect 257160 97854 257212 97860
rect 257172 95470 257200 97854
rect 257344 97300 257396 97306
rect 257344 97242 257396 97248
rect 257252 96960 257304 96966
rect 257252 96902 257304 96908
rect 257160 95464 257212 95470
rect 257160 95406 257212 95412
rect 257068 71052 257120 71058
rect 257068 70994 257120 71000
rect 256976 32428 257028 32434
rect 256976 32370 257028 32376
rect 257264 3262 257292 96902
rect 257356 95554 257384 97242
rect 257448 95690 257476 100028
rect 257632 97442 257660 100028
rect 257620 97436 257672 97442
rect 257620 97378 257672 97384
rect 257448 95662 257844 95690
rect 257356 95526 257476 95554
rect 257344 95464 257396 95470
rect 257344 95406 257396 95412
rect 257356 80782 257384 95406
rect 257448 93226 257476 95526
rect 257816 93854 257844 95662
rect 257908 94586 257936 100028
rect 257896 94580 257948 94586
rect 257896 94522 257948 94528
rect 257816 93826 258028 93854
rect 257436 93220 257488 93226
rect 257436 93162 257488 93168
rect 257344 80776 257396 80782
rect 257344 80718 257396 80724
rect 258000 21418 258028 93826
rect 258184 83570 258212 100028
rect 258382 100014 258488 100042
rect 258172 83564 258224 83570
rect 258172 83506 258224 83512
rect 258460 54602 258488 100014
rect 258644 97918 258672 100028
rect 258632 97912 258684 97918
rect 258632 97854 258684 97860
rect 258828 84194 258856 100028
rect 259104 84194 259132 100028
rect 259380 97782 259408 100028
rect 259578 100014 259684 100042
rect 259368 97776 259420 97782
rect 259368 97718 259420 97724
rect 258736 84166 258856 84194
rect 259012 84166 259132 84194
rect 258736 82210 258764 84166
rect 258724 82204 258776 82210
rect 258724 82146 258776 82152
rect 259012 58750 259040 84166
rect 259000 58744 259052 58750
rect 259000 58686 259052 58692
rect 259656 57322 259684 100014
rect 259644 57316 259696 57322
rect 259644 57258 259696 57264
rect 258448 54596 258500 54602
rect 258448 54538 258500 54544
rect 259840 38010 259868 100028
rect 260116 97016 260144 100028
rect 260300 97646 260328 100028
rect 260392 100014 260590 100042
rect 260288 97640 260340 97646
rect 260288 97582 260340 97588
rect 260024 96988 260144 97016
rect 259920 96960 259972 96966
rect 259920 96902 259972 96908
rect 259828 38004 259880 38010
rect 259828 37946 259880 37952
rect 259932 36650 259960 96902
rect 260024 75274 260052 96988
rect 260392 96966 260420 100014
rect 260380 96960 260432 96966
rect 260380 96902 260432 96908
rect 260104 96892 260156 96898
rect 260104 96834 260156 96840
rect 260012 75268 260064 75274
rect 260012 75210 260064 75216
rect 259920 36644 259972 36650
rect 259920 36586 259972 36592
rect 257988 21412 258040 21418
rect 257988 21354 258040 21360
rect 258080 19984 258132 19990
rect 258080 19926 258132 19932
rect 258092 16574 258120 19926
rect 258092 16546 258304 16574
rect 257252 3256 257304 3262
rect 257252 3198 257304 3204
rect 258276 480 258304 16546
rect 259460 10464 259512 10470
rect 259460 10406 259512 10412
rect 259472 3534 259500 10406
rect 260116 10402 260144 96834
rect 260196 96756 260248 96762
rect 260196 96698 260248 96704
rect 260208 86358 260236 96698
rect 260852 87718 260880 100028
rect 261036 96898 261064 100028
rect 261116 96960 261168 96966
rect 261116 96902 261168 96908
rect 261024 96892 261076 96898
rect 261024 96834 261076 96840
rect 260840 87712 260892 87718
rect 260840 87654 260892 87660
rect 260196 86352 260248 86358
rect 260196 86294 260248 86300
rect 261128 73914 261156 96902
rect 261312 84194 261340 100028
rect 261404 100014 261602 100042
rect 261404 96966 261432 100014
rect 261392 96960 261444 96966
rect 261392 96902 261444 96908
rect 261484 96892 261536 96898
rect 261484 96834 261536 96840
rect 261392 96824 261444 96830
rect 261392 96766 261444 96772
rect 261220 84166 261340 84194
rect 261116 73908 261168 73914
rect 261116 73850 261168 73856
rect 261220 35290 261248 84166
rect 261208 35284 261260 35290
rect 261208 35226 261260 35232
rect 260932 21412 260984 21418
rect 260932 21354 260984 21360
rect 260944 16574 260972 21354
rect 261404 20058 261432 96766
rect 261496 79490 261524 96834
rect 261772 84194 261800 100028
rect 261864 100014 262062 100042
rect 261864 96830 261892 100014
rect 261852 96824 261904 96830
rect 261852 96766 261904 96772
rect 262232 96762 262260 100028
rect 262220 96756 262272 96762
rect 262220 96698 262272 96704
rect 262508 89078 262536 100028
rect 262588 96960 262640 96966
rect 262588 96902 262640 96908
rect 262496 89072 262548 89078
rect 262496 89014 262548 89020
rect 261680 84166 261800 84194
rect 261484 79484 261536 79490
rect 261484 79426 261536 79432
rect 261680 55962 261708 84166
rect 261668 55956 261720 55962
rect 261668 55898 261720 55904
rect 262600 33862 262628 96902
rect 262784 84194 262812 100028
rect 262968 96898 262996 100028
rect 263060 100014 263258 100042
rect 263336 100014 263534 100042
rect 262956 96892 263008 96898
rect 262956 96834 263008 96840
rect 263060 90438 263088 100014
rect 263336 96966 263364 100014
rect 263324 96960 263376 96966
rect 263324 96902 263376 96908
rect 263048 90432 263100 90438
rect 263048 90374 263100 90380
rect 263704 84194 263732 100028
rect 263980 94586 264008 100028
rect 264072 100014 264270 100042
rect 263968 94580 264020 94586
rect 263968 94522 264020 94528
rect 264072 89714 264100 100014
rect 264440 99374 264468 100028
rect 264348 99346 264468 99374
rect 264532 100014 264730 100042
rect 264152 94784 264204 94790
rect 264152 94726 264204 94732
rect 262692 84166 262812 84194
rect 263612 84166 263732 84194
rect 263796 89686 264100 89714
rect 262692 60110 262720 84166
rect 263612 72554 263640 84166
rect 263600 72548 263652 72554
rect 263600 72490 263652 72496
rect 262680 60104 262732 60110
rect 262680 60046 262732 60052
rect 262588 33856 262640 33862
rect 262588 33798 262640 33804
rect 263796 31142 263824 89686
rect 264164 84194 264192 94726
rect 264348 89714 264376 99346
rect 264532 94790 264560 100014
rect 264520 94784 264572 94790
rect 264520 94726 264572 94732
rect 264520 94580 264572 94586
rect 264520 94522 264572 94528
rect 264348 89686 264468 89714
rect 264440 84194 264468 89686
rect 264072 84166 264192 84194
rect 264348 84166 264468 84194
rect 263784 31136 263836 31142
rect 263784 31078 263836 31084
rect 264072 21486 264100 84166
rect 264348 69766 264376 84166
rect 264336 69760 264388 69766
rect 264336 69702 264388 69708
rect 264532 24206 264560 94522
rect 264992 29714 265020 100028
rect 265176 97306 265204 100028
rect 265268 100014 265466 100042
rect 265544 100014 265742 100042
rect 265164 97300 265216 97306
rect 265164 97242 265216 97248
rect 265164 90160 265216 90166
rect 265164 90102 265216 90108
rect 265072 66904 265124 66910
rect 265072 66846 265124 66852
rect 264980 29708 265032 29714
rect 264980 29650 265032 29656
rect 264520 24200 264572 24206
rect 264520 24142 264572 24148
rect 264060 21480 264112 21486
rect 264060 21422 264112 21428
rect 261392 20052 261444 20058
rect 261392 19994 261444 20000
rect 260944 16546 261800 16574
rect 260104 10396 260156 10402
rect 260104 10338 260156 10344
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 260656 3528 260708 3534
rect 260656 3470 260708 3476
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 259472 480 259500 3334
rect 260668 480 260696 3470
rect 261772 480 261800 16546
rect 264152 11824 264204 11830
rect 264152 11766 264204 11772
rect 262956 3596 263008 3602
rect 262956 3538 263008 3544
rect 262968 480 262996 3538
rect 264164 480 264192 11766
rect 257038 354 257150 480
rect 256804 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265084 354 265112 66846
rect 265176 53174 265204 90102
rect 265268 68406 265296 100014
rect 265440 96756 265492 96762
rect 265440 96698 265492 96704
rect 265452 90506 265480 96698
rect 265440 90500 265492 90506
rect 265440 90442 265492 90448
rect 265544 90166 265572 100014
rect 265624 96688 265676 96694
rect 265624 96630 265676 96636
rect 265532 90160 265584 90166
rect 265532 90102 265584 90108
rect 265256 68400 265308 68406
rect 265256 68342 265308 68348
rect 265164 53168 265216 53174
rect 265164 53110 265216 53116
rect 265636 22846 265664 96630
rect 265912 91934 265940 100028
rect 265900 91928 265952 91934
rect 265900 91870 265952 91876
rect 266188 84194 266216 100028
rect 266386 100014 266492 100042
rect 266096 84166 266216 84194
rect 266096 67046 266124 84166
rect 266084 67040 266136 67046
rect 266084 66982 266136 66988
rect 266464 51814 266492 100014
rect 266648 97646 266676 100028
rect 266636 97640 266688 97646
rect 266636 97582 266688 97588
rect 266728 94580 266780 94586
rect 266728 94522 266780 94528
rect 266452 51808 266504 51814
rect 266452 51750 266504 51756
rect 266740 50454 266768 94522
rect 266924 89714 266952 100028
rect 267108 94586 267136 100028
rect 267384 96762 267412 100028
rect 267476 100014 267674 100042
rect 267372 96756 267424 96762
rect 267372 96698 267424 96704
rect 267096 94580 267148 94586
rect 267096 94522 267148 94528
rect 266832 89686 266952 89714
rect 266832 76702 266860 89686
rect 266820 76696 266872 76702
rect 266820 76638 266872 76644
rect 267476 65686 267504 100014
rect 267844 94518 267872 100028
rect 267924 94784 267976 94790
rect 267924 94726 267976 94732
rect 267832 94512 267884 94518
rect 267832 94454 267884 94460
rect 267740 87644 267792 87650
rect 267740 87586 267792 87592
rect 267464 65680 267516 65686
rect 267464 65622 267516 65628
rect 266728 50448 266780 50454
rect 266728 50390 266780 50396
rect 265624 22840 265676 22846
rect 265624 22782 265676 22788
rect 267752 3738 267780 87586
rect 267832 83496 267884 83502
rect 267832 83438 267884 83444
rect 267740 3732 267792 3738
rect 267740 3674 267792 3680
rect 266544 3664 266596 3670
rect 266544 3606 266596 3612
rect 266556 480 266584 3606
rect 267844 3482 267872 83438
rect 267936 47666 267964 94726
rect 268120 89146 268148 100028
rect 268292 97844 268344 97850
rect 268292 97786 268344 97792
rect 268200 94852 268252 94858
rect 268200 94794 268252 94800
rect 268108 89140 268160 89146
rect 268108 89082 268160 89088
rect 268212 87786 268240 94794
rect 268304 89714 268332 97786
rect 268396 96694 268424 100028
rect 268384 96688 268436 96694
rect 268384 96630 268436 96636
rect 268476 96688 268528 96694
rect 268476 96630 268528 96636
rect 268304 89686 268424 89714
rect 268200 87780 268252 87786
rect 268200 87722 268252 87728
rect 267924 47660 267976 47666
rect 267924 47602 267976 47608
rect 268396 6390 268424 89686
rect 268488 83638 268516 96630
rect 268580 94790 268608 100028
rect 268672 100014 268870 100042
rect 268672 94858 268700 100014
rect 268660 94852 268712 94858
rect 268660 94794 268712 94800
rect 268568 94784 268620 94790
rect 268568 94726 268620 94732
rect 269132 94586 269160 100028
rect 269330 100014 269436 100042
rect 269120 94580 269172 94586
rect 269120 94522 269172 94528
rect 268660 94512 268712 94518
rect 268660 94454 268712 94460
rect 268476 83632 268528 83638
rect 268476 83574 268528 83580
rect 268672 75342 268700 94454
rect 268660 75336 268712 75342
rect 268660 75278 268712 75284
rect 269408 73982 269436 100014
rect 269592 96082 269620 100028
rect 269776 99374 269804 100028
rect 269684 99346 269804 99374
rect 269868 100014 270066 100042
rect 269580 96076 269632 96082
rect 269580 96018 269632 96024
rect 269396 73976 269448 73982
rect 269396 73918 269448 73924
rect 269684 62966 269712 99346
rect 269764 97368 269816 97374
rect 269764 97310 269816 97316
rect 269672 62960 269724 62966
rect 269672 62902 269724 62908
rect 268384 6384 268436 6390
rect 268384 6326 268436 6332
rect 269776 4962 269804 97310
rect 269868 25634 269896 100014
rect 270132 94580 270184 94586
rect 270132 94522 270184 94528
rect 270144 64326 270172 94522
rect 270328 86426 270356 100028
rect 270526 100014 270632 100042
rect 270500 96892 270552 96898
rect 270500 96834 270552 96840
rect 270512 94654 270540 96834
rect 270500 94648 270552 94654
rect 270500 94590 270552 94596
rect 270604 94518 270632 100014
rect 270592 94512 270644 94518
rect 270592 94454 270644 94460
rect 270592 94376 270644 94382
rect 270592 94318 270644 94324
rect 270316 86420 270368 86426
rect 270316 86362 270368 86368
rect 270132 64320 270184 64326
rect 270132 64262 270184 64268
rect 270604 43518 270632 94318
rect 270788 84194 270816 100028
rect 271064 96694 271092 100028
rect 271052 96688 271104 96694
rect 271052 96630 271104 96636
rect 270868 94580 270920 94586
rect 270868 94522 270920 94528
rect 270696 84166 270816 84194
rect 270696 46374 270724 84166
rect 270880 82278 270908 94522
rect 270868 82272 270920 82278
rect 270868 82214 270920 82220
rect 270684 46368 270736 46374
rect 270684 46310 270736 46316
rect 270592 43512 270644 43518
rect 270592 43454 270644 43460
rect 269856 25628 269908 25634
rect 269856 25570 269908 25576
rect 270776 13252 270828 13258
rect 270776 13194 270828 13200
rect 269764 4956 269816 4962
rect 269764 4898 269816 4904
rect 268476 3732 268528 3738
rect 268476 3674 268528 3680
rect 270040 3732 270092 3738
rect 270040 3674 270092 3680
rect 267752 3454 267872 3482
rect 267752 480 267780 3454
rect 265318 354 265430 480
rect 265084 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 3674
rect 270052 480 270080 3674
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 13194
rect 271248 13190 271276 100028
rect 271328 94512 271380 94518
rect 271328 94454 271380 94460
rect 271340 61538 271368 94454
rect 271524 94382 271552 100028
rect 271616 100014 271814 100042
rect 271616 94586 271644 100014
rect 271604 94580 271656 94586
rect 271604 94522 271656 94528
rect 271512 94376 271564 94382
rect 271512 94318 271564 94324
rect 271984 93294 272012 100028
rect 272064 94580 272116 94586
rect 272064 94522 272116 94528
rect 271972 93288 272024 93294
rect 271972 93230 272024 93236
rect 272076 78130 272104 94522
rect 272260 84194 272288 100028
rect 272536 96898 272564 100028
rect 272524 96892 272576 96898
rect 272524 96834 272576 96840
rect 272720 94586 272748 100028
rect 272812 100014 273010 100042
rect 272708 94580 272760 94586
rect 272708 94522 272760 94528
rect 272168 84166 272288 84194
rect 272064 78124 272116 78130
rect 272064 78066 272116 78072
rect 271328 61532 271380 61538
rect 271328 61474 271380 61480
rect 272168 42226 272196 84166
rect 272812 72622 272840 100014
rect 273272 93362 273300 100028
rect 273260 93356 273312 93362
rect 273260 93298 273312 93304
rect 272800 72616 272852 72622
rect 272800 72558 272852 72564
rect 273456 71126 273484 100028
rect 273732 96218 273760 100028
rect 273916 96778 273944 100028
rect 273824 96750 273944 96778
rect 273996 96824 274048 96830
rect 273996 96766 274048 96772
rect 273720 96212 273772 96218
rect 273720 96154 273772 96160
rect 273824 84930 273852 96750
rect 273904 96688 273956 96694
rect 273904 96630 273956 96636
rect 273812 84924 273864 84930
rect 273812 84866 273864 84872
rect 273444 71120 273496 71126
rect 273444 71062 273496 71068
rect 272156 42220 272208 42226
rect 272156 42162 272208 42168
rect 271236 13184 271288 13190
rect 271236 13126 271288 13132
rect 273916 7818 273944 96630
rect 274008 60178 274036 96766
rect 274192 84194 274220 100028
rect 274100 84166 274220 84194
rect 274284 100014 274482 100042
rect 273996 60172 274048 60178
rect 273996 60114 274048 60120
rect 274100 15978 274128 84166
rect 274284 40866 274312 100014
rect 274364 97640 274416 97646
rect 274364 97582 274416 97588
rect 274376 96694 274404 97582
rect 274364 96688 274416 96694
rect 274364 96630 274416 96636
rect 274652 92002 274680 100028
rect 274928 96830 274956 100028
rect 275204 98002 275232 100028
rect 275112 97974 275232 98002
rect 275008 96892 275060 96898
rect 275008 96834 275060 96840
rect 274916 96824 274968 96830
rect 274916 96766 274968 96772
rect 274640 91996 274692 92002
rect 274640 91938 274692 91944
rect 274272 40860 274324 40866
rect 274272 40802 274324 40808
rect 275020 27062 275048 96834
rect 275112 69834 275140 97974
rect 275388 97900 275416 100028
rect 275204 97872 275416 97900
rect 275204 96354 275232 97872
rect 275376 97776 275428 97782
rect 275376 97718 275428 97724
rect 275284 97572 275336 97578
rect 275284 97514 275336 97520
rect 275192 96348 275244 96354
rect 275192 96290 275244 96296
rect 275100 69828 275152 69834
rect 275100 69770 275152 69776
rect 275008 27056 275060 27062
rect 275008 26998 275060 27004
rect 274088 15972 274140 15978
rect 274088 15914 274140 15920
rect 273904 7812 273956 7818
rect 273904 7754 273956 7760
rect 275296 5030 275324 97514
rect 275388 49162 275416 97718
rect 275468 96960 275520 96966
rect 275468 96902 275520 96908
rect 275480 90574 275508 96902
rect 275468 90568 275520 90574
rect 275468 90510 275520 90516
rect 275664 84194 275692 100028
rect 275756 100014 275954 100042
rect 275756 96898 275784 100014
rect 276124 96966 276152 100028
rect 276112 96960 276164 96966
rect 276112 96902 276164 96908
rect 276204 96960 276256 96966
rect 276204 96902 276256 96908
rect 275744 96892 275796 96898
rect 275744 96834 275796 96840
rect 276216 86494 276244 96902
rect 276400 92070 276428 100028
rect 276492 100014 276690 100042
rect 276388 92064 276440 92070
rect 276388 92006 276440 92012
rect 276204 86488 276256 86494
rect 276204 86430 276256 86436
rect 275572 84166 275692 84194
rect 275572 80850 275600 84166
rect 275560 80844 275612 80850
rect 275560 80786 275612 80792
rect 276492 68474 276520 100014
rect 276860 97986 276888 100028
rect 276952 100014 277150 100042
rect 276848 97980 276900 97986
rect 276848 97922 276900 97928
rect 276664 97436 276716 97442
rect 276664 97378 276716 97384
rect 276480 68468 276532 68474
rect 276480 68410 276532 68416
rect 275376 49156 275428 49162
rect 275376 49098 275428 49104
rect 276676 39506 276704 97378
rect 276952 84998 276980 100014
rect 277320 96966 277348 100028
rect 277610 100014 277716 100042
rect 277308 96960 277360 96966
rect 277308 96902 277360 96908
rect 277688 89214 277716 100014
rect 277676 89208 277728 89214
rect 277676 89150 277728 89156
rect 276940 84992 276992 84998
rect 276940 84934 276992 84940
rect 277872 84194 277900 100028
rect 278056 97442 278084 100028
rect 278044 97436 278096 97442
rect 278044 97378 278096 97384
rect 278044 97028 278096 97034
rect 278044 96970 278096 96976
rect 277780 84166 277900 84194
rect 277780 58818 277808 84166
rect 277768 58812 277820 58818
rect 277768 58754 277820 58760
rect 276664 39500 276716 39506
rect 276664 39442 276716 39448
rect 277952 14544 278004 14550
rect 277952 14486 278004 14492
rect 276020 6384 276072 6390
rect 276020 6326 276072 6332
rect 275284 5024 275336 5030
rect 275284 4966 275336 4972
rect 272432 4956 272484 4962
rect 272432 4898 272484 4904
rect 272444 480 272472 4898
rect 274824 4344 274876 4350
rect 274824 4286 274876 4292
rect 273628 3800 273680 3806
rect 273628 3742 273680 3748
rect 273640 480 273668 3742
rect 274836 480 274864 4286
rect 276032 480 276060 6326
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 277136 480 277164 3810
rect 277964 3482 277992 14486
rect 278056 4894 278084 96970
rect 278136 96688 278188 96694
rect 278136 96630 278188 96636
rect 278148 6254 278176 96630
rect 278332 84194 278360 100028
rect 278240 84166 278360 84194
rect 278424 100014 278622 100042
rect 278806 100014 278912 100042
rect 278240 79558 278268 84166
rect 278228 79552 278280 79558
rect 278228 79494 278280 79500
rect 278424 17406 278452 100014
rect 278884 44946 278912 100014
rect 279068 94722 279096 100028
rect 279344 97782 279372 100028
rect 279542 100014 279648 100042
rect 279332 97776 279384 97782
rect 279332 97718 279384 97724
rect 279424 97436 279476 97442
rect 279424 97378 279476 97384
rect 279148 97096 279200 97102
rect 279148 97038 279200 97044
rect 279056 94716 279108 94722
rect 279056 94658 279108 94664
rect 278872 44940 278924 44946
rect 278872 44882 278924 44888
rect 278412 17400 278464 17406
rect 278412 17342 278464 17348
rect 279160 7614 279188 97038
rect 279148 7608 279200 7614
rect 279148 7550 279200 7556
rect 278136 6248 278188 6254
rect 278136 6190 278188 6196
rect 278044 4888 278096 4894
rect 278044 4830 278096 4836
rect 279436 4350 279464 97378
rect 279620 96966 279648 100014
rect 279608 96960 279660 96966
rect 279608 96902 279660 96908
rect 279516 96892 279568 96898
rect 279516 96834 279568 96840
rect 279528 10334 279556 96834
rect 279804 84194 279832 100028
rect 279896 100014 280094 100042
rect 279896 97102 279924 100014
rect 279884 97096 279936 97102
rect 279884 97038 279936 97044
rect 279884 96960 279936 96966
rect 279884 96902 279936 96908
rect 279896 87854 279924 96902
rect 280264 96898 280292 100028
rect 280540 97034 280568 100028
rect 280816 97374 280844 100028
rect 280804 97368 280856 97374
rect 280804 97310 280856 97316
rect 280528 97028 280580 97034
rect 280528 96970 280580 96976
rect 281000 96948 281028 100028
rect 281276 97850 281304 100028
rect 281264 97844 281316 97850
rect 281264 97786 281316 97792
rect 280632 96920 281028 96948
rect 280252 96892 280304 96898
rect 280252 96834 280304 96840
rect 279884 87848 279936 87854
rect 279884 87790 279936 87796
rect 279712 84166 279832 84194
rect 279712 76770 279740 84166
rect 279700 76764 279752 76770
rect 279700 76706 279752 76712
rect 279516 10328 279568 10334
rect 279516 10270 279568 10276
rect 280632 9042 280660 96920
rect 280804 96824 280856 96830
rect 280804 96766 280856 96772
rect 280816 9110 280844 96766
rect 281460 96694 281488 100028
rect 281736 97646 281764 100028
rect 281724 97640 281776 97646
rect 281724 97582 281776 97588
rect 281816 96960 281868 96966
rect 281816 96902 281868 96908
rect 281448 96688 281500 96694
rect 281448 96630 281500 96636
rect 281828 18630 281856 96902
rect 282012 84194 282040 100028
rect 282196 96966 282224 100028
rect 282288 100014 282486 100042
rect 282564 100014 282762 100042
rect 282946 100014 283052 100042
rect 282184 96960 282236 96966
rect 282184 96902 282236 96908
rect 282184 96756 282236 96762
rect 282184 96698 282236 96704
rect 281920 84166 282040 84194
rect 281816 18624 281868 18630
rect 281816 18566 281868 18572
rect 280804 9104 280856 9110
rect 280804 9046 280856 9052
rect 280620 9036 280672 9042
rect 280620 8978 280672 8984
rect 281920 7750 281948 84166
rect 281908 7744 281960 7750
rect 281908 7686 281960 7692
rect 281908 6928 281960 6934
rect 281908 6870 281960 6876
rect 279424 4344 279476 4350
rect 279424 4286 279476 4292
rect 279516 3936 279568 3942
rect 279516 3878 279568 3884
rect 277964 3454 278360 3482
rect 278332 480 278360 3454
rect 279528 480 279556 3878
rect 280712 3324 280764 3330
rect 280712 3266 280764 3272
rect 280724 480 280752 3266
rect 281920 480 281948 6870
rect 282196 6186 282224 96698
rect 282184 6180 282236 6186
rect 282184 6122 282236 6128
rect 282288 4826 282316 100014
rect 282564 8974 282592 100014
rect 283024 11762 283052 100014
rect 283208 96762 283236 100028
rect 283484 97578 283512 100028
rect 283472 97572 283524 97578
rect 283472 97514 283524 97520
rect 283288 96960 283340 96966
rect 283288 96902 283340 96908
rect 283196 96756 283248 96762
rect 283196 96698 283248 96704
rect 283012 11756 283064 11762
rect 283012 11698 283064 11704
rect 282552 8968 282604 8974
rect 282552 8910 282604 8916
rect 283300 6322 283328 96902
rect 283668 84194 283696 100028
rect 283944 84194 283972 100028
rect 284036 100014 284234 100042
rect 284036 96966 284064 100014
rect 284024 96960 284076 96966
rect 284024 96902 284076 96908
rect 284404 96830 284432 100028
rect 284680 96966 284708 100028
rect 284668 96960 284720 96966
rect 284668 96902 284720 96908
rect 284392 96824 284444 96830
rect 284392 96766 284444 96772
rect 284484 95396 284536 95402
rect 284484 95338 284536 95344
rect 283576 84166 283696 84194
rect 283852 84166 283972 84194
rect 283576 14482 283604 84166
rect 283564 14476 283616 14482
rect 283564 14418 283616 14424
rect 283852 13122 283880 84166
rect 283840 13116 283892 13122
rect 283840 13058 283892 13064
rect 284496 10470 284524 95338
rect 284864 84194 284892 100028
rect 284944 97980 284996 97986
rect 284944 97922 284996 97928
rect 284772 84166 284892 84194
rect 284772 80714 284800 84166
rect 284760 80708 284812 80714
rect 284760 80650 284812 80656
rect 284484 10464 284536 10470
rect 284484 10406 284536 10412
rect 284956 6390 284984 97922
rect 285140 84194 285168 100028
rect 285220 96960 285272 96966
rect 285220 96902 285272 96908
rect 285048 84166 285168 84194
rect 285048 19990 285076 84166
rect 285036 19984 285088 19990
rect 285036 19926 285088 19932
rect 284944 6384 284996 6390
rect 284944 6326 284996 6332
rect 283288 6316 283340 6322
rect 283288 6258 283340 6264
rect 282276 4820 282328 4826
rect 282276 4762 282328 4768
rect 284300 4140 284352 4146
rect 284300 4082 284352 4088
rect 283104 4072 283156 4078
rect 283104 4014 283156 4020
rect 283116 480 283144 4014
rect 284312 480 284340 4082
rect 285232 3466 285260 96902
rect 285416 84194 285444 100028
rect 285600 95402 285628 100028
rect 285588 95396 285640 95402
rect 285588 95338 285640 95344
rect 285324 84166 285444 84194
rect 285220 3460 285272 3466
rect 285220 3402 285272 3408
rect 285324 3398 285352 84166
rect 285692 3602 285720 100098
rect 285890 100014 285996 100042
rect 285968 21418 285996 100014
rect 286336 84194 286364 100028
rect 286416 96960 286468 96966
rect 286416 96902 286468 96908
rect 286244 84166 286364 84194
rect 285956 21412 286008 21418
rect 285956 21354 286008 21360
rect 286244 11830 286272 84166
rect 286232 11824 286284 11830
rect 286232 11766 286284 11772
rect 286428 3670 286456 96902
rect 286612 93922 286640 100028
rect 286704 100014 286902 100042
rect 287086 100014 287192 100042
rect 286704 96966 286732 100014
rect 287164 96966 287192 100014
rect 287348 97186 287376 100028
rect 287256 97158 287376 97186
rect 287440 100014 287638 100042
rect 286692 96960 286744 96966
rect 286692 96902 286744 96908
rect 287152 96960 287204 96966
rect 287152 96902 287204 96908
rect 287256 96898 287284 97158
rect 287440 97050 287468 100014
rect 287348 97022 287468 97050
rect 287244 96892 287296 96898
rect 287244 96834 287296 96840
rect 287348 96778 287376 97022
rect 287428 96960 287480 96966
rect 287428 96902 287480 96908
rect 286520 93894 286640 93922
rect 287164 96750 287376 96778
rect 286520 66910 286548 93894
rect 286508 66904 286560 66910
rect 286508 66846 286560 66852
rect 287164 3738 287192 96750
rect 287244 96688 287296 96694
rect 287244 96630 287296 96636
rect 287256 87650 287284 96630
rect 287244 87644 287296 87650
rect 287244 87586 287296 87592
rect 287440 83502 287468 96902
rect 287808 84194 287836 100028
rect 287888 96960 287940 96966
rect 287888 96902 287940 96908
rect 287716 84166 287836 84194
rect 287428 83496 287480 83502
rect 287428 83438 287480 83444
rect 287716 13258 287744 84166
rect 287704 13252 287756 13258
rect 287704 13194 287756 13200
rect 287900 3806 287928 96902
rect 288084 93922 288112 100028
rect 288176 100014 288374 100042
rect 288176 96966 288204 100014
rect 288544 97442 288572 100028
rect 288820 97986 288848 100028
rect 288808 97980 288860 97986
rect 288808 97922 288860 97928
rect 288532 97436 288584 97442
rect 288532 97378 288584 97384
rect 288164 96960 288216 96966
rect 288164 96902 288216 96908
rect 287992 93894 288112 93922
rect 287992 4962 288020 93894
rect 289004 84194 289032 100028
rect 289084 96892 289136 96898
rect 289084 96834 289136 96840
rect 288636 84166 289032 84194
rect 287980 4956 288032 4962
rect 287980 4898 288032 4904
rect 288636 3874 288664 84166
rect 289096 6934 289124 96834
rect 289280 84194 289308 100028
rect 289188 84166 289308 84194
rect 289372 100014 289570 100042
rect 289188 14550 289216 84166
rect 289176 14544 289228 14550
rect 289176 14486 289228 14492
rect 289084 6928 289136 6934
rect 289084 6870 289136 6876
rect 289372 3942 289400 100014
rect 289740 84194 289768 100028
rect 290016 96898 290044 100028
rect 290096 96960 290148 96966
rect 290096 96902 290148 96908
rect 290004 96892 290056 96898
rect 290004 96834 290056 96840
rect 289648 84166 289768 84194
rect 289360 3936 289412 3942
rect 289360 3878 289412 3884
rect 288624 3868 288676 3874
rect 288624 3810 288676 3816
rect 287888 3800 287940 3806
rect 287888 3742 287940 3748
rect 287152 3732 287204 3738
rect 287152 3674 287204 3680
rect 286416 3664 286468 3670
rect 286416 3606 286468 3612
rect 285680 3596 285732 3602
rect 285680 3538 285732 3544
rect 286600 3596 286652 3602
rect 286600 3538 286652 3544
rect 285404 3528 285456 3534
rect 285404 3470 285456 3476
rect 285312 3392 285364 3398
rect 285312 3334 285364 3340
rect 285416 480 285444 3470
rect 286612 480 286640 3538
rect 289648 3330 289676 84166
rect 290108 3602 290136 96902
rect 290292 84194 290320 100028
rect 290476 84194 290504 100028
rect 290200 84166 290320 84194
rect 290384 84166 290504 84194
rect 290568 100014 290766 100042
rect 290844 100014 291042 100042
rect 290200 4078 290228 84166
rect 290384 4146 290412 84166
rect 290372 4140 290424 4146
rect 290372 4082 290424 4088
rect 290188 4072 290240 4078
rect 290188 4014 290240 4020
rect 290096 3596 290148 3602
rect 290096 3538 290148 3544
rect 290568 3534 290596 100014
rect 290844 96966 290872 100014
rect 290832 96960 290884 96966
rect 290832 96902 290884 96908
rect 290556 3528 290608 3534
rect 290556 3470 290608 3476
rect 289636 3324 289688 3330
rect 289636 3266 289688 3272
rect 290188 3324 290240 3330
rect 290188 3266 290240 3272
rect 288992 3188 289044 3194
rect 288992 3130 289044 3136
rect 287796 3120 287848 3126
rect 287796 3062 287848 3068
rect 287808 480 287836 3062
rect 289004 480 289032 3130
rect 290200 480 290228 3266
rect 291212 3126 291240 100028
rect 291304 100014 291502 100042
rect 291304 3194 291332 100014
rect 291568 96960 291620 96966
rect 291568 96902 291620 96908
rect 291580 3602 291608 96902
rect 291764 84194 291792 100028
rect 291948 84194 291976 100028
rect 291672 84166 291792 84194
rect 291856 84166 291976 84194
rect 292040 100014 292238 100042
rect 291568 3596 291620 3602
rect 291568 3538 291620 3544
rect 291672 3330 291700 84166
rect 291660 3324 291712 3330
rect 291660 3266 291712 3272
rect 291292 3188 291344 3194
rect 291292 3130 291344 3136
rect 291200 3120 291252 3126
rect 291200 3062 291252 3068
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 354 291466 480
rect 291856 354 291884 84166
rect 292040 3466 292068 100014
rect 292408 96966 292436 100028
rect 292396 96960 292448 96966
rect 292396 96902 292448 96908
rect 292684 84194 292712 100028
rect 292764 96960 292816 96966
rect 292764 96902 292816 96908
rect 292592 84166 292712 84194
rect 292592 16574 292620 84166
rect 292592 16546 292712 16574
rect 292684 4146 292712 16546
rect 292672 4140 292724 4146
rect 292672 4082 292724 4088
rect 292776 4010 292804 96902
rect 292960 84194 292988 100028
rect 293144 96966 293172 100028
rect 293236 100014 293434 100042
rect 293512 100014 293710 100042
rect 293132 96960 293184 96966
rect 293132 96902 293184 96908
rect 292868 84166 292988 84194
rect 292868 4078 292896 84166
rect 292856 4072 292908 4078
rect 292856 4014 292908 4020
rect 292764 4004 292816 4010
rect 292764 3946 292816 3952
rect 293236 3942 293264 100014
rect 293512 5506 293540 100014
rect 293880 84194 293908 100028
rect 293788 84166 293908 84194
rect 293972 100014 294170 100042
rect 293788 9110 293816 84166
rect 293776 9104 293828 9110
rect 293776 9046 293828 9052
rect 293500 5500 293552 5506
rect 293500 5442 293552 5448
rect 293224 3936 293276 3942
rect 293224 3878 293276 3884
rect 293972 3874 294000 100014
rect 294432 97646 294460 100028
rect 294420 97640 294472 97646
rect 294420 97582 294472 97588
rect 294236 96960 294288 96966
rect 294236 96902 294288 96908
rect 293960 3868 294012 3874
rect 293960 3810 294012 3816
rect 293684 3596 293736 3602
rect 293684 3538 293736 3544
rect 292028 3460 292080 3466
rect 292028 3402 292080 3408
rect 292580 3460 292632 3466
rect 292580 3402 292632 3408
rect 292592 480 292620 3402
rect 293696 480 293724 3538
rect 294248 3398 294276 96902
rect 294616 84862 294644 100028
rect 294708 100014 294906 100042
rect 294984 100014 295182 100042
rect 294708 96966 294736 100014
rect 294696 96960 294748 96966
rect 294696 96902 294748 96908
rect 294604 84856 294656 84862
rect 294604 84798 294656 84804
rect 294984 84194 295012 100014
rect 295352 97510 295380 100028
rect 295628 97578 295656 100028
rect 295616 97572 295668 97578
rect 295616 97514 295668 97520
rect 295340 97504 295392 97510
rect 295340 97446 295392 97452
rect 295432 97096 295484 97102
rect 295432 97038 295484 97044
rect 294708 84166 295012 84194
rect 294708 10402 294736 84166
rect 294696 10396 294748 10402
rect 294696 10338 294748 10344
rect 295444 4894 295472 97038
rect 295812 84194 295840 100028
rect 295904 100014 296102 100042
rect 296180 100014 296378 100042
rect 295904 97102 295932 100014
rect 295892 97096 295944 97102
rect 295892 97038 295944 97044
rect 295892 96960 295944 96966
rect 295892 96902 295944 96908
rect 295720 84166 295840 84194
rect 295720 4962 295748 84166
rect 295904 6118 295932 96902
rect 296180 7682 296208 100014
rect 296548 96966 296576 100028
rect 296536 96960 296588 96966
rect 296536 96902 296588 96908
rect 296824 84194 296852 100028
rect 296904 97096 296956 97102
rect 296904 97038 296956 97044
rect 296732 84166 296852 84194
rect 296732 66910 296760 84166
rect 296720 66904 296772 66910
rect 296720 66846 296772 66852
rect 296168 7676 296220 7682
rect 296168 7618 296220 7624
rect 296916 6322 296944 97038
rect 297100 84194 297128 100028
rect 297284 97442 297312 100028
rect 297376 100014 297574 100042
rect 297652 100014 297850 100042
rect 297272 97436 297324 97442
rect 297272 97378 297324 97384
rect 297376 97102 297404 100014
rect 297364 97096 297416 97102
rect 297364 97038 297416 97044
rect 297364 96960 297416 96966
rect 297364 96902 297416 96908
rect 297008 84166 297128 84194
rect 297008 18630 297036 84166
rect 296996 18624 297048 18630
rect 296996 18566 297048 18572
rect 297376 7614 297404 96902
rect 297652 20126 297680 100014
rect 298020 96966 298048 100028
rect 298296 97034 298324 100028
rect 298284 97028 298336 97034
rect 298284 96970 298336 96976
rect 298008 96960 298060 96966
rect 298008 96902 298060 96908
rect 298376 96960 298428 96966
rect 298376 96902 298428 96908
rect 298100 96892 298152 96898
rect 298100 96834 298152 96840
rect 297640 20120 297692 20126
rect 297640 20062 297692 20068
rect 298112 9042 298140 96834
rect 298388 14618 298416 96902
rect 298572 84194 298600 100028
rect 298756 97306 298784 100028
rect 298848 100014 299046 100042
rect 299124 100014 299322 100042
rect 298744 97300 298796 97306
rect 298744 97242 298796 97248
rect 298848 96966 298876 100014
rect 298836 96960 298888 96966
rect 298836 96902 298888 96908
rect 299124 96898 299152 100014
rect 299112 96892 299164 96898
rect 299112 96834 299164 96840
rect 298480 84166 298600 84194
rect 298480 58682 298508 84166
rect 298468 58676 298520 58682
rect 298468 58618 298520 58624
rect 298376 14612 298428 14618
rect 298376 14554 298428 14560
rect 298100 9036 298152 9042
rect 298100 8978 298152 8984
rect 299492 8974 299520 100028
rect 299572 96960 299624 96966
rect 299572 96902 299624 96908
rect 299480 8968 299532 8974
rect 299480 8910 299532 8916
rect 297364 7608 297416 7614
rect 297364 7550 297416 7556
rect 296904 6316 296956 6322
rect 296904 6258 296956 6264
rect 295892 6112 295944 6118
rect 295892 6054 295944 6060
rect 295708 4956 295760 4962
rect 295708 4898 295760 4904
rect 295432 4888 295484 4894
rect 295432 4830 295484 4836
rect 299584 4826 299612 96902
rect 299768 84194 299796 100028
rect 299952 96966 299980 100028
rect 299940 96960 299992 96966
rect 299940 96902 299992 96908
rect 300032 96960 300084 96966
rect 300032 96902 300084 96908
rect 299676 84166 299796 84194
rect 299676 15910 299704 84166
rect 300044 26926 300072 96902
rect 300228 95946 300256 100028
rect 300320 100014 300518 100042
rect 300216 95940 300268 95946
rect 300216 95882 300268 95888
rect 300320 53106 300348 100014
rect 300688 96966 300716 100028
rect 300964 97374 300992 100028
rect 300952 97368 301004 97374
rect 300952 97310 301004 97316
rect 301044 97096 301096 97102
rect 301044 97038 301096 97044
rect 300676 96960 300728 96966
rect 300676 96902 300728 96908
rect 300308 53100 300360 53106
rect 300308 53042 300360 53048
rect 300032 26920 300084 26926
rect 300032 26862 300084 26868
rect 299664 15904 299716 15910
rect 299664 15846 299716 15852
rect 301056 11762 301084 97038
rect 301240 84194 301268 100028
rect 301424 84194 301452 100028
rect 301516 100014 301714 100042
rect 301792 100014 301990 100042
rect 301516 97102 301544 100014
rect 301504 97096 301556 97102
rect 301504 97038 301556 97044
rect 301792 96948 301820 100014
rect 301148 84166 301268 84194
rect 301332 84166 301452 84194
rect 301516 96920 301820 96948
rect 301148 60178 301176 84166
rect 301136 60172 301188 60178
rect 301136 60114 301188 60120
rect 301332 42090 301360 84166
rect 301320 42084 301372 42090
rect 301320 42026 301372 42032
rect 301516 17270 301544 96920
rect 302160 84194 302188 100028
rect 302240 97640 302292 97646
rect 302240 97582 302292 97588
rect 301792 84166 302188 84194
rect 301792 29646 301820 84166
rect 301780 29640 301832 29646
rect 301780 29582 301832 29588
rect 301504 17264 301556 17270
rect 301504 17206 301556 17212
rect 301044 11756 301096 11762
rect 301044 11698 301096 11704
rect 300768 9104 300820 9110
rect 300768 9046 300820 9052
rect 299664 5500 299716 5506
rect 299664 5442 299716 5448
rect 299572 4820 299624 4826
rect 299572 4762 299624 4768
rect 294880 4140 294932 4146
rect 294880 4082 294932 4088
rect 294236 3392 294288 3398
rect 294236 3334 294288 3340
rect 294892 480 294920 4082
rect 296076 4072 296128 4078
rect 296076 4014 296128 4020
rect 296088 480 296116 4014
rect 297272 4004 297324 4010
rect 297272 3946 297324 3952
rect 297284 480 297312 3946
rect 298468 3936 298520 3942
rect 298468 3878 298520 3884
rect 298480 480 298508 3878
rect 299676 480 299704 5442
rect 300780 480 300808 9046
rect 302252 6914 302280 97582
rect 302436 84194 302464 100028
rect 302516 96960 302568 96966
rect 302516 96902 302568 96908
rect 302344 84166 302464 84194
rect 302344 82142 302372 84166
rect 302332 82136 302384 82142
rect 302332 82078 302384 82084
rect 302528 13122 302556 96902
rect 302712 84194 302740 100028
rect 302896 84194 302924 100028
rect 302988 100014 303186 100042
rect 302988 96966 303016 100014
rect 302976 96960 303028 96966
rect 302976 96902 303028 96908
rect 303356 84194 303384 100028
rect 303646 100014 303752 100042
rect 303724 97238 303752 100014
rect 303712 97232 303764 97238
rect 303712 97174 303764 97180
rect 303712 97096 303764 97102
rect 303712 97038 303764 97044
rect 303620 84856 303672 84862
rect 303620 84798 303672 84804
rect 302620 84166 302740 84194
rect 302804 84166 302924 84194
rect 302988 84166 303384 84194
rect 302620 69698 302648 84166
rect 302608 69692 302660 69698
rect 302608 69634 302660 69640
rect 302804 39506 302832 84166
rect 302792 39500 302844 39506
rect 302792 39442 302844 39448
rect 302988 28286 303016 84166
rect 302976 28280 303028 28286
rect 302976 28222 303028 28228
rect 302516 13116 302568 13122
rect 302516 13058 302568 13064
rect 302252 6886 303200 6914
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 301976 480 302004 3810
rect 303172 480 303200 6886
rect 291354 326 291884 354
rect 291354 -960 291466 326
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303632 354 303660 84798
rect 303724 6254 303752 97038
rect 303908 84194 303936 100028
rect 304092 84194 304120 100028
rect 304184 100014 304382 100042
rect 304184 97102 304212 100014
rect 304448 97232 304500 97238
rect 304448 97174 304500 97180
rect 304172 97096 304224 97102
rect 304172 97038 304224 97044
rect 304172 96960 304224 96966
rect 304172 96902 304224 96908
rect 303816 84166 303936 84194
rect 304000 84166 304120 84194
rect 303816 71058 303844 84166
rect 303804 71052 303856 71058
rect 303804 70994 303856 71000
rect 304000 46306 304028 84166
rect 303988 46300 304040 46306
rect 303988 46242 304040 46248
rect 304184 32502 304212 96902
rect 304460 75410 304488 97174
rect 304644 93430 304672 100028
rect 304828 96966 304856 100028
rect 304816 96960 304868 96966
rect 304816 96902 304868 96908
rect 304632 93424 304684 93430
rect 304632 93366 304684 93372
rect 305104 84194 305132 100028
rect 305184 97096 305236 97102
rect 305184 97038 305236 97044
rect 305012 84166 305132 84194
rect 304448 75404 304500 75410
rect 304448 75346 304500 75352
rect 304172 32496 304224 32502
rect 304172 32438 304224 32444
rect 305012 31210 305040 84166
rect 305000 31204 305052 31210
rect 305000 31146 305052 31152
rect 305196 14482 305224 97038
rect 305380 94790 305408 100028
rect 305368 94784 305420 94790
rect 305368 94726 305420 94732
rect 305564 84194 305592 100028
rect 305656 100014 305854 100042
rect 305932 100014 306130 100042
rect 305656 97102 305684 100014
rect 305644 97096 305696 97102
rect 305644 97038 305696 97044
rect 305736 97028 305788 97034
rect 305736 96970 305788 96976
rect 305644 96960 305696 96966
rect 305644 96902 305696 96908
rect 305472 84166 305592 84194
rect 305472 74050 305500 84166
rect 305460 74044 305512 74050
rect 305460 73986 305512 73992
rect 305656 72622 305684 96902
rect 305644 72616 305696 72622
rect 305644 72558 305696 72564
rect 305184 14476 305236 14482
rect 305184 14418 305236 14424
rect 305748 10334 305776 96970
rect 305932 92002 305960 100014
rect 306300 96966 306328 100028
rect 306288 96960 306340 96966
rect 306288 96902 306340 96908
rect 306380 96892 306432 96898
rect 306380 96834 306432 96840
rect 305920 91996 305972 92002
rect 305920 91938 305972 91944
rect 306392 20058 306420 96834
rect 306576 84194 306604 100028
rect 306656 96960 306708 96966
rect 306656 96902 306708 96908
rect 306668 86426 306696 96902
rect 306852 90574 306880 100028
rect 307036 97594 307064 100028
rect 306944 97566 307064 97594
rect 307128 100014 307326 100042
rect 306944 94722 306972 97566
rect 307024 97504 307076 97510
rect 307024 97446 307076 97452
rect 306932 94716 306984 94722
rect 306932 94658 306984 94664
rect 306840 90568 306892 90574
rect 306840 90510 306892 90516
rect 306656 86420 306708 86426
rect 306656 86362 306708 86368
rect 306484 84166 306604 84194
rect 306484 61538 306512 84166
rect 306472 61532 306524 61538
rect 306472 61474 306524 61480
rect 306380 20052 306432 20058
rect 306380 19994 306432 20000
rect 306380 10396 306432 10402
rect 306380 10338 306432 10344
rect 305736 10328 305788 10334
rect 305736 10270 305788 10276
rect 303712 6248 303764 6254
rect 303712 6190 303764 6196
rect 305552 3392 305604 3398
rect 305552 3334 305604 3340
rect 305564 480 305592 3334
rect 304326 354 304438 480
rect 303632 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 10338
rect 307036 4214 307064 97446
rect 307128 96898 307156 100014
rect 307208 97572 307260 97578
rect 307208 97514 307260 97520
rect 307116 96892 307168 96898
rect 307116 96834 307168 96840
rect 307220 84194 307248 97514
rect 307496 96966 307524 100028
rect 307484 96960 307536 96966
rect 307484 96902 307536 96908
rect 307772 96218 307800 100028
rect 307852 96960 307904 96966
rect 307852 96902 307904 96908
rect 307760 96212 307812 96218
rect 307760 96154 307812 96160
rect 307128 84166 307248 84194
rect 307128 8294 307156 84166
rect 307864 62966 307892 96902
rect 308048 85066 308076 100028
rect 308232 96830 308260 100028
rect 308324 100014 308522 100042
rect 308600 100014 308798 100042
rect 308220 96824 308272 96830
rect 308220 96766 308272 96772
rect 308036 85060 308088 85066
rect 308036 85002 308088 85008
rect 308324 80918 308352 100014
rect 308600 96966 308628 100014
rect 308588 96960 308640 96966
rect 308588 96902 308640 96908
rect 308968 96150 308996 100028
rect 308956 96144 309008 96150
rect 308956 96086 309008 96092
rect 309244 84194 309272 100028
rect 309324 96960 309376 96966
rect 309324 96902 309376 96908
rect 309152 84166 309272 84194
rect 308312 80912 308364 80918
rect 308312 80854 308364 80860
rect 309152 69834 309180 84166
rect 309140 69828 309192 69834
rect 309140 69770 309192 69776
rect 307852 62960 307904 62966
rect 307852 62902 307904 62908
rect 309336 11830 309364 96902
rect 309520 84194 309548 100028
rect 309704 87854 309732 100028
rect 309796 100014 309994 100042
rect 310072 100014 310270 100042
rect 309692 87848 309744 87854
rect 309692 87790 309744 87796
rect 309428 84166 309548 84194
rect 309428 13258 309456 84166
rect 309796 73982 309824 100014
rect 310072 96966 310100 100014
rect 310060 96960 310112 96966
rect 310060 96902 310112 96908
rect 310440 84194 310468 100028
rect 310520 96960 310572 96966
rect 310520 96902 310572 96908
rect 310072 84166 310468 84194
rect 310072 83706 310100 84166
rect 310060 83700 310112 83706
rect 310060 83642 310112 83648
rect 309784 73976 309836 73982
rect 309784 73918 309836 73924
rect 310532 26994 310560 96902
rect 310716 93922 310744 100028
rect 310900 96966 310928 100028
rect 311176 97594 311204 100028
rect 311084 97566 311204 97594
rect 311268 100014 311466 100042
rect 310888 96960 310940 96966
rect 310888 96902 310940 96908
rect 310980 95396 311032 95402
rect 310980 95338 311032 95344
rect 310624 93894 310744 93922
rect 310624 71194 310652 93894
rect 310992 72554 311020 95338
rect 311084 84998 311112 97566
rect 311164 97436 311216 97442
rect 311164 97378 311216 97384
rect 311072 84992 311124 84998
rect 311072 84934 311124 84940
rect 310980 72548 311032 72554
rect 310980 72490 311032 72496
rect 310612 71188 310664 71194
rect 310612 71130 310664 71136
rect 310520 26988 310572 26994
rect 310520 26930 310572 26936
rect 309416 13252 309468 13258
rect 309416 13194 309468 13200
rect 309324 11824 309376 11830
rect 309324 11766 309376 11772
rect 307116 8288 307168 8294
rect 307116 8230 307168 8236
rect 309048 8288 309100 8294
rect 309048 8230 309100 8236
rect 307024 4208 307076 4214
rect 307024 4150 307076 4156
rect 307944 4208 307996 4214
rect 307944 4150 307996 4156
rect 307956 480 307984 4150
rect 309060 480 309088 8230
rect 310244 4956 310296 4962
rect 310244 4898 310296 4904
rect 310256 480 310284 4898
rect 311176 4486 311204 97378
rect 311268 95402 311296 100014
rect 311256 95396 311308 95402
rect 311256 95338 311308 95344
rect 311636 94654 311664 100028
rect 311912 97578 311940 100028
rect 311900 97572 311952 97578
rect 311900 97514 311952 97520
rect 311992 96892 312044 96898
rect 311992 96834 312044 96840
rect 311624 94648 311676 94654
rect 311624 94590 311676 94596
rect 312004 17338 312032 96834
rect 312188 84194 312216 100028
rect 312372 84194 312400 100028
rect 312452 96960 312504 96966
rect 312452 96902 312504 96908
rect 312096 84166 312216 84194
rect 312280 84166 312400 84194
rect 312096 82278 312124 84166
rect 312084 82272 312136 82278
rect 312084 82214 312136 82220
rect 312280 75342 312308 84166
rect 312464 79490 312492 96902
rect 312648 91934 312676 100028
rect 312740 100014 312938 100042
rect 312740 96966 312768 100014
rect 312728 96960 312780 96966
rect 312728 96902 312780 96908
rect 313108 96898 313136 100028
rect 313096 96892 313148 96898
rect 313096 96834 313148 96840
rect 312636 91928 312688 91934
rect 312636 91870 312688 91876
rect 313384 90506 313412 100028
rect 313464 96960 313516 96966
rect 313464 96902 313516 96908
rect 313372 90500 313424 90506
rect 313372 90442 313424 90448
rect 312452 79484 312504 79490
rect 312452 79426 312504 79432
rect 312268 75336 312320 75342
rect 312268 75278 312320 75284
rect 311992 17332 312044 17338
rect 311992 17274 312044 17280
rect 312636 7676 312688 7682
rect 312636 7618 312688 7624
rect 311440 4888 311492 4894
rect 311440 4830 311492 4836
rect 311164 4480 311216 4486
rect 311164 4422 311216 4428
rect 311452 480 311480 4830
rect 312648 480 312676 7618
rect 313476 6186 313504 96902
rect 313660 93922 313688 100028
rect 313844 96966 313872 100028
rect 313832 96960 313884 96966
rect 313832 96902 313884 96908
rect 313924 96960 313976 96966
rect 313924 96902 313976 96908
rect 313568 93894 313688 93922
rect 313568 60110 313596 93894
rect 313556 60104 313608 60110
rect 313556 60046 313608 60052
rect 313936 25634 313964 96902
rect 314120 84194 314148 100028
rect 314212 100014 314410 100042
rect 314212 96966 314240 100014
rect 314200 96960 314252 96966
rect 314200 96902 314252 96908
rect 314580 84194 314608 100028
rect 314660 96960 314712 96966
rect 314660 96902 314712 96908
rect 314028 84166 314148 84194
rect 314212 84166 314608 84194
rect 314028 80850 314056 84166
rect 314016 80844 314068 80850
rect 314016 80786 314068 80792
rect 314212 32434 314240 84166
rect 314200 32428 314252 32434
rect 314200 32370 314252 32376
rect 313924 25628 313976 25634
rect 313924 25570 313976 25576
rect 314672 24206 314700 96902
rect 314856 84194 314884 100028
rect 315040 84194 315068 100028
rect 314764 84166 314884 84194
rect 314948 84166 315068 84194
rect 315132 100014 315330 100042
rect 315408 100014 315606 100042
rect 314764 68474 314792 84166
rect 314752 68468 314804 68474
rect 314752 68410 314804 68416
rect 314752 66904 314804 66910
rect 314752 66846 314804 66852
rect 314660 24200 314712 24206
rect 314660 24142 314712 24148
rect 313464 6180 313516 6186
rect 313464 6122 313516 6128
rect 313832 6112 313884 6118
rect 313832 6054 313884 6060
rect 313844 480 313872 6054
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314764 354 314792 66846
rect 314948 57390 314976 84166
rect 314936 57384 314988 57390
rect 314936 57326 314988 57332
rect 315132 29714 315160 100014
rect 315304 96824 315356 96830
rect 315304 96766 315356 96772
rect 315316 89214 315344 96766
rect 315304 89208 315356 89214
rect 315304 89150 315356 89156
rect 315408 67046 315436 100014
rect 315776 96966 315804 100028
rect 315764 96960 315816 96966
rect 315764 96902 315816 96908
rect 315396 67040 315448 67046
rect 315396 66982 315448 66988
rect 316052 64326 316080 100028
rect 316132 96960 316184 96966
rect 316132 96902 316184 96908
rect 316040 64320 316092 64326
rect 316040 64262 316092 64268
rect 315120 29708 315172 29714
rect 315120 29650 315172 29656
rect 316144 28354 316172 96902
rect 316328 96830 316356 100028
rect 316316 96824 316368 96830
rect 316316 96766 316368 96772
rect 316512 86290 316540 100028
rect 316604 100014 316802 100042
rect 316604 96966 316632 100014
rect 317064 97646 317092 100028
rect 317052 97640 317104 97646
rect 317052 97582 317104 97588
rect 316592 96960 316644 96966
rect 316592 96902 316644 96908
rect 316500 86284 316552 86290
rect 316500 86226 316552 86232
rect 317248 84194 317276 100028
rect 317524 84194 317552 100028
rect 317604 96960 317656 96966
rect 317604 96902 317656 96908
rect 316604 84166 317276 84194
rect 317432 84166 317552 84194
rect 316604 78130 316632 84166
rect 316592 78124 316644 78130
rect 316592 78066 316644 78072
rect 316132 28348 316184 28354
rect 316132 28290 316184 28296
rect 316040 18624 316092 18630
rect 316040 18566 316092 18572
rect 316052 16574 316080 18566
rect 316052 16546 316264 16574
rect 316236 480 316264 16546
rect 317432 14550 317460 84166
rect 317616 22846 317644 96902
rect 317800 84194 317828 100028
rect 317984 84194 318012 100028
rect 317708 84166 317828 84194
rect 317892 84166 318012 84194
rect 318076 100014 318274 100042
rect 317708 79422 317736 84166
rect 317696 79416 317748 79422
rect 317696 79358 317748 79364
rect 317892 56030 317920 84166
rect 317880 56024 317932 56030
rect 317880 55966 317932 55972
rect 318076 31142 318104 100014
rect 318444 84194 318472 100028
rect 318536 100014 318734 100042
rect 318536 96966 318564 100014
rect 318524 96960 318576 96966
rect 318524 96902 318576 96908
rect 318800 96960 318852 96966
rect 318800 96902 318852 96908
rect 318352 84166 318472 84194
rect 318352 65686 318380 84166
rect 318340 65680 318392 65686
rect 318340 65622 318392 65628
rect 318064 31136 318116 31142
rect 318064 31078 318116 31084
rect 317604 22840 317656 22846
rect 317604 22782 317656 22788
rect 318812 19990 318840 96902
rect 318996 84194 319024 100028
rect 319180 89146 319208 100028
rect 319272 100014 319470 100042
rect 319548 100014 319746 100042
rect 319168 89140 319220 89146
rect 319168 89082 319220 89088
rect 318904 84166 319024 84194
rect 318904 60042 318932 84166
rect 318892 60036 318944 60042
rect 318892 59978 318944 59984
rect 319272 21486 319300 100014
rect 319444 97300 319496 97306
rect 319444 97242 319496 97248
rect 319260 21480 319312 21486
rect 319260 21422 319312 21428
rect 318892 20120 318944 20126
rect 318892 20062 318944 20068
rect 318800 19984 318852 19990
rect 318800 19926 318852 19932
rect 318904 16574 318932 20062
rect 318904 16546 319392 16574
rect 317420 14544 317472 14550
rect 317420 14486 317472 14492
rect 318524 6316 318576 6322
rect 318524 6258 318576 6264
rect 317328 4480 317380 4486
rect 317328 4422 317380 4428
rect 317340 480 317368 4422
rect 318536 480 318564 6258
rect 319364 3482 319392 16546
rect 319456 4214 319484 97242
rect 319548 96966 319576 100014
rect 319536 96960 319588 96966
rect 319536 96902 319588 96908
rect 319916 84194 319944 100028
rect 319548 84166 319944 84194
rect 319548 64258 319576 84166
rect 319536 64252 319588 64258
rect 319536 64194 319588 64200
rect 320192 54670 320220 100028
rect 320284 100014 320482 100042
rect 320180 54664 320232 54670
rect 320180 54606 320232 54612
rect 320284 13190 320312 100014
rect 320652 84194 320680 100028
rect 320560 84166 320680 84194
rect 320744 100014 320942 100042
rect 320560 78062 320588 84166
rect 320548 78056 320600 78062
rect 320548 77998 320600 78004
rect 320744 18698 320772 100014
rect 321204 96082 321232 100028
rect 321192 96076 321244 96082
rect 321192 96018 321244 96024
rect 321388 84194 321416 100028
rect 321664 84194 321692 100028
rect 321744 96960 321796 96966
rect 321744 96902 321796 96908
rect 321020 84166 321416 84194
rect 321572 84166 321692 84194
rect 321020 62898 321048 84166
rect 321572 69766 321600 84166
rect 321560 69760 321612 69766
rect 321560 69702 321612 69708
rect 321008 62892 321060 62898
rect 321008 62834 321060 62840
rect 320732 18692 320784 18698
rect 320732 18634 320784 18640
rect 320272 13184 320324 13190
rect 320272 13126 320324 13132
rect 321652 10328 321704 10334
rect 321652 10270 321704 10276
rect 320916 7608 320968 7614
rect 320916 7550 320968 7556
rect 319444 4208 319496 4214
rect 319444 4150 319496 4156
rect 319364 3454 319760 3482
rect 319732 480 319760 3454
rect 320928 480 320956 7550
rect 321664 3482 321692 10270
rect 321756 3602 321784 96902
rect 321940 84194 321968 100028
rect 322124 97782 322152 100028
rect 322216 100014 322414 100042
rect 322112 97776 322164 97782
rect 322112 97718 322164 97724
rect 321848 84166 321968 84194
rect 321848 58818 321876 84166
rect 321836 58812 321888 58818
rect 321836 58754 321888 58760
rect 322216 51814 322244 100014
rect 322584 96966 322612 100028
rect 322676 100014 322874 100042
rect 322572 96960 322624 96966
rect 322572 96902 322624 96908
rect 322676 87786 322704 100014
rect 322940 96960 322992 96966
rect 322940 96902 322992 96908
rect 322664 87780 322716 87786
rect 322664 87722 322716 87728
rect 322204 51808 322256 51814
rect 322204 51750 322256 51756
rect 321744 3596 321796 3602
rect 321744 3538 321796 3544
rect 321664 3454 322152 3482
rect 322124 480 322152 3454
rect 322952 3330 322980 96902
rect 323136 84194 323164 100028
rect 323320 96966 323348 100028
rect 323308 96960 323360 96966
rect 323308 96902 323360 96908
rect 323400 96960 323452 96966
rect 323596 96948 323624 100028
rect 323400 96902 323452 96908
rect 323504 96920 323624 96948
rect 323688 100014 323886 100042
rect 323044 84166 323164 84194
rect 323044 73914 323072 84166
rect 323032 73908 323084 73914
rect 323032 73850 323084 73856
rect 323032 58676 323084 58682
rect 323032 58618 323084 58624
rect 322940 3324 322992 3330
rect 322940 3266 322992 3272
rect 314998 354 315110 480
rect 314764 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323044 354 323072 58618
rect 323412 3398 323440 96902
rect 323504 58750 323532 96920
rect 323584 96824 323636 96830
rect 323584 96766 323636 96772
rect 323596 86358 323624 96766
rect 323584 86352 323636 86358
rect 323584 86294 323636 86300
rect 323492 58744 323544 58750
rect 323492 58686 323544 58692
rect 323688 50454 323716 100014
rect 324056 96966 324084 100028
rect 324044 96960 324096 96966
rect 324044 96902 324096 96908
rect 324332 76702 324360 100028
rect 324412 96960 324464 96966
rect 324412 96902 324464 96908
rect 324320 76696 324372 76702
rect 324320 76638 324372 76644
rect 323676 50448 323728 50454
rect 323676 50390 323728 50396
rect 324320 4208 324372 4214
rect 324320 4150 324372 4156
rect 324332 3482 324360 4150
rect 324424 4078 324452 96902
rect 324608 84194 324636 100028
rect 324792 84194 324820 100028
rect 324516 84166 324636 84194
rect 324700 84166 324820 84194
rect 324884 100014 325082 100042
rect 325160 100014 325358 100042
rect 324516 53174 324544 84166
rect 324504 53168 324556 53174
rect 324504 53110 324556 53116
rect 324596 14612 324648 14618
rect 324596 14554 324648 14560
rect 324412 4072 324464 4078
rect 324412 4014 324464 4020
rect 324608 3482 324636 14554
rect 324700 4146 324728 84166
rect 324884 57322 324912 100014
rect 325160 89078 325188 100014
rect 325528 96966 325556 100028
rect 325804 97034 325832 100028
rect 325792 97028 325844 97034
rect 325792 96970 325844 96976
rect 325516 96960 325568 96966
rect 325516 96902 325568 96908
rect 325148 89072 325200 89078
rect 325148 89014 325200 89020
rect 325988 84194 326016 100028
rect 325896 84166 326016 84194
rect 326080 100014 326278 100042
rect 325896 71126 325924 84166
rect 325884 71120 325936 71126
rect 325884 71062 325936 71068
rect 324872 57316 324924 57322
rect 324872 57258 324924 57264
rect 324688 4140 324740 4146
rect 324688 4082 324740 4088
rect 326080 4010 326108 100014
rect 326344 95804 326396 95810
rect 326344 95746 326396 95752
rect 326068 4004 326120 4010
rect 326068 3946 326120 3952
rect 326356 3942 326384 95746
rect 326540 93294 326568 100028
rect 326528 93288 326580 93294
rect 326528 93230 326580 93236
rect 326724 84194 326752 100028
rect 326816 100014 327014 100042
rect 326816 95810 326844 100014
rect 327080 97096 327132 97102
rect 327080 97038 327132 97044
rect 326804 95804 326856 95810
rect 326804 95746 326856 95752
rect 326632 84166 326752 84194
rect 326632 80782 326660 84166
rect 326620 80776 326672 80782
rect 326620 80718 326672 80724
rect 326804 9036 326856 9042
rect 326804 8978 326856 8984
rect 326344 3936 326396 3942
rect 326344 3878 326396 3884
rect 324332 3454 324452 3482
rect 324608 3454 325648 3482
rect 323400 3392 323452 3398
rect 323400 3334 323452 3340
rect 324424 480 324452 3454
rect 325620 480 325648 3454
rect 326816 480 326844 8978
rect 327092 3874 327120 97038
rect 327276 84194 327304 100028
rect 327460 84194 327488 100028
rect 327552 100014 327750 100042
rect 327828 100014 328026 100042
rect 327552 97102 327580 100014
rect 327540 97096 327592 97102
rect 327540 97038 327592 97044
rect 327724 97028 327776 97034
rect 327724 96970 327776 96976
rect 327540 96960 327592 96966
rect 327540 96902 327592 96908
rect 327184 84166 327304 84194
rect 327368 84166 327488 84194
rect 327184 55962 327212 84166
rect 327172 55956 327224 55962
rect 327172 55898 327224 55904
rect 327368 25566 327396 84166
rect 327356 25560 327408 25566
rect 327356 25502 327408 25508
rect 327552 24138 327580 96902
rect 327736 83570 327764 96970
rect 327724 83564 327776 83570
rect 327724 83506 327776 83512
rect 327828 54602 327856 100014
rect 328196 96966 328224 100028
rect 328184 96960 328236 96966
rect 328184 96902 328236 96908
rect 327816 54596 327868 54602
rect 327816 54538 327868 54544
rect 327540 24132 327592 24138
rect 327540 24074 327592 24080
rect 328000 8968 328052 8974
rect 328000 8910 328052 8916
rect 327080 3868 327132 3874
rect 327080 3810 327132 3816
rect 328012 480 328040 8910
rect 328472 3806 328500 100028
rect 328552 97096 328604 97102
rect 328552 97038 328604 97044
rect 328460 3800 328512 3806
rect 328460 3742 328512 3748
rect 328564 3738 328592 97038
rect 328748 97034 328776 100028
rect 328736 97028 328788 97034
rect 328736 96970 328788 96976
rect 328932 84194 328960 100028
rect 329024 100014 329222 100042
rect 329300 100014 329498 100042
rect 329024 97102 329052 100014
rect 329012 97096 329064 97102
rect 329012 97038 329064 97044
rect 329012 96960 329064 96966
rect 329012 96902 329064 96908
rect 328840 84166 328960 84194
rect 328840 72486 328868 84166
rect 328828 72480 328880 72486
rect 328828 72422 328880 72428
rect 329024 22778 329052 96902
rect 329300 51746 329328 100014
rect 329668 96966 329696 100028
rect 329656 96960 329708 96966
rect 329656 96902 329708 96908
rect 329944 84194 329972 100028
rect 330128 96830 330156 100028
rect 330208 96960 330260 96966
rect 330208 96902 330260 96908
rect 330116 96824 330168 96830
rect 330116 96766 330168 96772
rect 329852 84166 329972 84194
rect 329288 51740 329340 51746
rect 329288 51682 329340 51688
rect 329012 22772 329064 22778
rect 329012 22714 329064 22720
rect 328736 15904 328788 15910
rect 328736 15846 328788 15852
rect 328552 3732 328604 3738
rect 328552 3674 328604 3680
rect 323278 354 323390 480
rect 323044 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 15846
rect 329852 3670 329880 84166
rect 329840 3664 329892 3670
rect 329840 3606 329892 3612
rect 330220 3534 330248 96902
rect 330404 87718 330432 100028
rect 330496 100014 330694 100042
rect 330496 96966 330524 100014
rect 330864 97510 330892 100028
rect 330956 100014 331154 100042
rect 330852 97504 330904 97510
rect 330852 97446 330904 97452
rect 330484 96960 330536 96966
rect 330484 96902 330536 96908
rect 330392 87712 330444 87718
rect 330392 87654 330444 87660
rect 330956 84194 330984 100014
rect 331220 95940 331272 95946
rect 331220 95882 331272 95888
rect 330496 84166 330984 84194
rect 330496 75274 330524 84166
rect 330484 75268 330536 75274
rect 330484 75210 330536 75216
rect 330392 4820 330444 4826
rect 330392 4762 330444 4768
rect 330208 3528 330260 3534
rect 330208 3470 330260 3476
rect 330404 480 330432 4762
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 95882
rect 331416 84194 331444 100028
rect 331600 97442 331628 100028
rect 331692 100014 331890 100042
rect 331968 100014 332166 100042
rect 331588 97436 331640 97442
rect 331588 97378 331640 97384
rect 331324 84166 331444 84194
rect 331324 49094 331352 84166
rect 331692 50386 331720 100014
rect 331864 97368 331916 97374
rect 331864 97310 331916 97316
rect 331680 50380 331732 50386
rect 331680 50322 331732 50328
rect 331312 49088 331364 49094
rect 331312 49030 331364 49036
rect 331876 4214 331904 97310
rect 331968 76634 331996 100014
rect 332140 97572 332192 97578
rect 332140 97514 332192 97520
rect 332048 96824 332100 96830
rect 332048 96766 332100 96772
rect 331956 76628 332008 76634
rect 331956 76570 332008 76576
rect 332060 68406 332088 96766
rect 332152 93362 332180 97514
rect 332336 97306 332364 100028
rect 332324 97300 332376 97306
rect 332324 97242 332376 97248
rect 332140 93356 332192 93362
rect 332140 93298 332192 93304
rect 332048 68400 332100 68406
rect 332048 68342 332100 68348
rect 332612 66978 332640 100028
rect 332692 96960 332744 96966
rect 332692 96902 332744 96908
rect 332600 66972 332652 66978
rect 332600 66914 332652 66920
rect 332600 53100 332652 53106
rect 332600 53042 332652 53048
rect 332612 16574 332640 53042
rect 332704 18630 332732 96902
rect 332888 84194 332916 100028
rect 333072 96014 333100 100028
rect 333164 100014 333362 100042
rect 333060 96008 333112 96014
rect 333060 95950 333112 95956
rect 332796 84166 332916 84194
rect 332796 21418 332824 84166
rect 333164 49026 333192 100014
rect 333336 97640 333388 97646
rect 333336 97582 333388 97588
rect 333244 97028 333296 97034
rect 333244 96970 333296 96976
rect 333256 53106 333284 96970
rect 333348 82210 333376 97582
rect 333532 96966 333560 100028
rect 333520 96960 333572 96966
rect 333520 96902 333572 96908
rect 333808 94586 333836 100028
rect 333796 94580 333848 94586
rect 333796 94522 333848 94528
rect 334084 84194 334112 100028
rect 334268 84194 334296 100028
rect 334544 97986 334572 100028
rect 334636 100014 334834 100042
rect 334532 97980 334584 97986
rect 334532 97922 334584 97928
rect 334348 96960 334400 96966
rect 334348 96902 334400 96908
rect 333992 84166 334112 84194
rect 334176 84166 334296 84194
rect 333336 82204 333388 82210
rect 333336 82146 333388 82152
rect 333992 65618 334020 84166
rect 333980 65612 334032 65618
rect 333980 65554 334032 65560
rect 333244 53100 333296 53106
rect 333244 53042 333296 53048
rect 333152 49020 333204 49026
rect 333152 48962 333204 48968
rect 332876 26920 332928 26926
rect 332876 26862 332928 26868
rect 332784 21412 332836 21418
rect 332784 21354 332836 21360
rect 332692 18624 332744 18630
rect 332692 18566 332744 18572
rect 332888 16574 332916 26862
rect 332612 16546 332732 16574
rect 332888 16546 333928 16574
rect 331864 4208 331916 4214
rect 331864 4150 331916 4156
rect 332704 480 332732 16546
rect 333900 480 333928 16546
rect 334176 4894 334204 84166
rect 334360 46238 334388 96902
rect 334636 47666 334664 100014
rect 335004 96966 335032 100028
rect 335280 97374 335308 100028
rect 335268 97368 335320 97374
rect 335268 97310 335320 97316
rect 334992 96960 335044 96966
rect 334992 96902 335044 96908
rect 335360 96960 335412 96966
rect 335360 96902 335412 96908
rect 334624 47660 334676 47666
rect 334624 47602 334676 47608
rect 334348 46232 334400 46238
rect 334348 46174 334400 46180
rect 335372 7614 335400 96902
rect 335452 60172 335504 60178
rect 335452 60114 335504 60120
rect 335464 16574 335492 60114
rect 335556 44946 335584 100028
rect 335636 97776 335688 97782
rect 335636 97718 335688 97724
rect 335648 96830 335676 97718
rect 335636 96824 335688 96830
rect 335636 96766 335688 96772
rect 335740 84194 335768 100028
rect 336016 97866 336044 100028
rect 335924 97838 336044 97866
rect 336108 100014 336306 100042
rect 335924 97646 335952 97838
rect 335912 97640 335964 97646
rect 335912 97582 335964 97588
rect 336108 97050 336136 100014
rect 336188 97980 336240 97986
rect 336188 97922 336240 97928
rect 335648 84166 335768 84194
rect 335832 97022 336136 97050
rect 335648 68338 335676 84166
rect 335636 68332 335688 68338
rect 335636 68274 335688 68280
rect 335544 44940 335596 44946
rect 335544 44882 335596 44888
rect 335832 43518 335860 97022
rect 336004 96824 336056 96830
rect 336004 96766 336056 96772
rect 336016 61470 336044 96766
rect 336200 93226 336228 97922
rect 336476 96966 336504 100028
rect 336464 96960 336516 96966
rect 336464 96902 336516 96908
rect 336188 93220 336240 93226
rect 336188 93162 336240 93168
rect 336752 91866 336780 100028
rect 336832 96892 336884 96898
rect 336832 96834 336884 96840
rect 336740 91860 336792 91866
rect 336740 91802 336792 91808
rect 336004 61464 336056 61470
rect 336004 61406 336056 61412
rect 335820 43512 335872 43518
rect 335820 43454 335872 43460
rect 336740 42084 336792 42090
rect 336740 42026 336792 42032
rect 335464 16546 336320 16574
rect 335360 7608 335412 7614
rect 335360 7550 335412 7556
rect 334164 4888 334216 4894
rect 334164 4830 334216 4836
rect 335084 4208 335136 4214
rect 335084 4150 335136 4156
rect 335096 480 335124 4150
rect 336292 480 336320 16546
rect 336752 6914 336780 42026
rect 336844 8974 336872 96834
rect 337028 84194 337056 100028
rect 337212 84194 337240 100028
rect 337292 96960 337344 96966
rect 337292 96902 337344 96908
rect 336936 84166 337056 84194
rect 337120 84166 337240 84194
rect 336936 42158 336964 84166
rect 337120 47598 337148 84166
rect 337108 47592 337160 47598
rect 337108 47534 337160 47540
rect 336924 42152 336976 42158
rect 336924 42094 336976 42100
rect 337304 40798 337332 96902
rect 337488 90438 337516 100028
rect 337672 96966 337700 100028
rect 337764 100014 337962 100042
rect 337660 96960 337712 96966
rect 337660 96902 337712 96908
rect 337764 96898 337792 100014
rect 338224 97578 338252 100028
rect 338212 97572 338264 97578
rect 338212 97514 338264 97520
rect 337752 96892 337804 96898
rect 337752 96834 337804 96840
rect 337476 90432 337528 90438
rect 337476 90374 337528 90380
rect 338408 84194 338436 100028
rect 338488 96892 338540 96898
rect 338488 96834 338540 96840
rect 338316 84166 338436 84194
rect 337292 40792 337344 40798
rect 337292 40734 337344 40740
rect 338316 39438 338344 84166
rect 338304 39432 338356 39438
rect 338304 39374 338356 39380
rect 338500 38010 338528 96834
rect 338684 84194 338712 100028
rect 338764 96960 338816 96966
rect 338764 96902 338816 96908
rect 338592 84166 338712 84194
rect 338592 57254 338620 84166
rect 338580 57248 338632 57254
rect 338580 57190 338632 57196
rect 338776 44878 338804 96902
rect 338960 89010 338988 100028
rect 339144 96898 339172 100028
rect 339236 100014 339434 100042
rect 339236 96966 339264 100014
rect 339224 96960 339276 96966
rect 339224 96902 339276 96908
rect 339500 96960 339552 96966
rect 339500 96902 339552 96908
rect 339132 96892 339184 96898
rect 339132 96834 339184 96840
rect 338948 89004 339000 89010
rect 338948 88946 339000 88952
rect 338764 44872 338816 44878
rect 338764 44814 338816 44820
rect 338488 38004 338540 38010
rect 338488 37946 338540 37952
rect 339512 15978 339540 96902
rect 339696 87650 339724 100028
rect 339880 96966 339908 100028
rect 339868 96960 339920 96966
rect 339868 96902 339920 96908
rect 339960 96960 340012 96966
rect 339960 96902 340012 96908
rect 339684 87644 339736 87650
rect 339684 87586 339736 87592
rect 339972 36650 340000 96902
rect 340156 84194 340184 100028
rect 340248 100014 340446 100042
rect 340248 84930 340276 100014
rect 340616 96966 340644 100028
rect 340604 96960 340656 96966
rect 340604 96902 340656 96908
rect 340892 96694 340920 100028
rect 340880 96688 340932 96694
rect 340880 96630 340932 96636
rect 340236 84924 340288 84930
rect 340236 84866 340288 84872
rect 341076 84194 341104 100028
rect 341156 96960 341208 96966
rect 341156 96902 341208 96908
rect 340064 84166 340184 84194
rect 340984 84166 341104 84194
rect 340064 43450 340092 84166
rect 340984 82142 341012 84166
rect 340880 82136 340932 82142
rect 340880 82078 340932 82084
rect 340972 82136 341024 82142
rect 340972 82078 341024 82084
rect 340052 43444 340104 43450
rect 340052 43386 340104 43392
rect 339960 36644 340012 36650
rect 339960 36586 340012 36592
rect 339592 17264 339644 17270
rect 339592 17206 339644 17212
rect 339500 15972 339552 15978
rect 339500 15914 339552 15920
rect 338672 11756 338724 11762
rect 338672 11698 338724 11704
rect 336832 8968 336884 8974
rect 336832 8910 336884 8916
rect 336752 6886 337056 6914
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 6886
rect 338684 480 338712 11698
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339604 354 339632 17206
rect 340892 2786 340920 82078
rect 340972 29640 341024 29646
rect 340972 29582 341024 29588
rect 340880 2780 340932 2786
rect 340880 2722 340932 2728
rect 340984 480 341012 29582
rect 341168 10334 341196 96902
rect 341352 84194 341380 100028
rect 341444 100014 341642 100042
rect 341444 96966 341472 100014
rect 341812 97850 341840 100028
rect 341904 100014 342102 100042
rect 341800 97844 341852 97850
rect 341800 97786 341852 97792
rect 341432 96960 341484 96966
rect 341432 96902 341484 96908
rect 341904 96778 341932 100014
rect 341260 84166 341380 84194
rect 341444 96750 341932 96778
rect 341260 64190 341288 84166
rect 341248 64184 341300 64190
rect 341248 64126 341300 64132
rect 341444 35290 341472 96750
rect 341892 96688 341944 96694
rect 341892 96630 341944 96636
rect 341904 42090 341932 96630
rect 342260 69692 342312 69698
rect 342260 69634 342312 69640
rect 341892 42084 341944 42090
rect 341892 42026 341944 42032
rect 341432 35284 341484 35290
rect 341432 35226 341484 35232
rect 342272 16574 342300 69634
rect 342364 66910 342392 100028
rect 342548 84194 342576 100028
rect 342628 96960 342680 96966
rect 342628 96902 342680 96908
rect 342456 84166 342576 84194
rect 342456 80714 342484 84166
rect 342444 80708 342496 80714
rect 342444 80650 342496 80656
rect 342352 66904 342404 66910
rect 342352 66846 342404 66852
rect 342640 31074 342668 96902
rect 342824 84194 342852 100028
rect 342732 84166 342852 84194
rect 342916 100014 343114 100042
rect 342732 33862 342760 84166
rect 342916 40730 342944 100014
rect 343284 84194 343312 100028
rect 343376 100014 343574 100042
rect 343376 96966 343404 100014
rect 343364 96960 343416 96966
rect 343364 96902 343416 96908
rect 343640 96892 343692 96898
rect 343640 96834 343692 96840
rect 343192 84166 343312 84194
rect 343192 79354 343220 84166
rect 343180 79348 343232 79354
rect 343180 79290 343232 79296
rect 342904 40724 342956 40730
rect 342904 40666 342956 40672
rect 343652 39370 343680 96834
rect 343836 84194 343864 100028
rect 344020 95946 344048 100028
rect 344100 96960 344152 96966
rect 344100 96902 344152 96908
rect 344008 95940 344060 95946
rect 344008 95882 344060 95888
rect 343744 84166 343864 84194
rect 343744 55894 343772 84166
rect 344112 77994 344140 96902
rect 344296 91798 344324 100028
rect 344388 100014 344586 100042
rect 344388 96898 344416 100014
rect 344756 96966 344784 100028
rect 344744 96960 344796 96966
rect 344744 96902 344796 96908
rect 344376 96892 344428 96898
rect 344376 96834 344428 96840
rect 344284 91792 344336 91798
rect 344284 91734 344336 91740
rect 344100 77988 344152 77994
rect 344100 77930 344152 77936
rect 343732 55888 343784 55894
rect 343732 55830 343784 55836
rect 343732 39500 343784 39506
rect 343732 39442 343784 39448
rect 343640 39364 343692 39370
rect 343640 39306 343692 39312
rect 342720 33856 342772 33862
rect 342720 33798 342772 33804
rect 342628 31068 342680 31074
rect 342628 31010 342680 31016
rect 343744 16574 343772 39442
rect 345032 29646 345060 100028
rect 345216 84194 345244 100028
rect 345492 97714 345520 100028
rect 345584 100014 345782 100042
rect 345480 97708 345532 97714
rect 345480 97650 345532 97656
rect 345296 96960 345348 96966
rect 345296 96902 345348 96908
rect 345124 84166 345244 84194
rect 345124 37942 345152 84166
rect 345112 37936 345164 37942
rect 345112 37878 345164 37884
rect 345308 36582 345336 96902
rect 345584 62830 345612 100014
rect 345952 96966 345980 100028
rect 346044 100014 346242 100042
rect 345940 96960 345992 96966
rect 345940 96902 345992 96908
rect 346044 76566 346072 100014
rect 346504 84194 346532 100028
rect 346688 84194 346716 100028
rect 346768 96960 346820 96966
rect 346768 96902 346820 96908
rect 346412 84166 346532 84194
rect 346596 84166 346716 84194
rect 346032 76560 346084 76566
rect 346032 76502 346084 76508
rect 345572 62824 345624 62830
rect 345572 62766 345624 62772
rect 346412 61402 346440 84166
rect 346400 61396 346452 61402
rect 346400 61338 346452 61344
rect 345296 36576 345348 36582
rect 345296 36518 345348 36524
rect 346596 35222 346624 84166
rect 346584 35216 346636 35222
rect 346584 35158 346636 35164
rect 345020 29640 345072 29646
rect 345020 29582 345072 29588
rect 346400 28280 346452 28286
rect 346400 28222 346452 28228
rect 342272 16546 342944 16574
rect 343744 16546 344600 16574
rect 341156 10328 341208 10334
rect 341156 10270 341208 10276
rect 342168 2780 342220 2786
rect 342168 2722 342220 2728
rect 342180 480 342208 2722
rect 339838 354 339950 480
rect 339604 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 345296 13116 345348 13122
rect 345296 13058 345348 13064
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 13058
rect 346412 6914 346440 28222
rect 346780 15910 346808 96902
rect 346964 94518 346992 100028
rect 347056 100014 347254 100042
rect 346952 94512 347004 94518
rect 346952 94454 347004 94460
rect 347056 28286 347084 100014
rect 347424 96966 347452 100028
rect 347516 100014 347714 100042
rect 347412 96960 347464 96966
rect 347412 96902 347464 96908
rect 347516 75206 347544 100014
rect 347780 96960 347832 96966
rect 347780 96902 347832 96908
rect 347792 84862 347820 96902
rect 347976 90370 348004 100028
rect 347964 90364 348016 90370
rect 347964 90306 348016 90312
rect 347780 84856 347832 84862
rect 347780 84798 347832 84804
rect 348160 84194 348188 100028
rect 348436 97034 348464 100028
rect 348424 97028 348476 97034
rect 348424 96970 348476 96976
rect 348620 96966 348648 100028
rect 348712 100014 348910 100042
rect 348608 96960 348660 96966
rect 348608 96902 348660 96908
rect 348712 84194 348740 100014
rect 349172 97782 349200 100028
rect 349160 97776 349212 97782
rect 349160 97718 349212 97724
rect 349356 84194 349384 100028
rect 349436 96892 349488 96898
rect 349436 96834 349488 96840
rect 348068 84166 348188 84194
rect 348252 84166 348740 84194
rect 349264 84166 349384 84194
rect 347780 75404 347832 75410
rect 347780 75346 347832 75352
rect 347504 75200 347556 75206
rect 347504 75142 347556 75148
rect 347044 28280 347096 28286
rect 347044 28222 347096 28228
rect 347792 16574 347820 75346
rect 348068 65550 348096 84166
rect 348056 65544 348108 65550
rect 348056 65486 348108 65492
rect 348252 33794 348280 84166
rect 349160 71052 349212 71058
rect 349160 70994 349212 71000
rect 348240 33788 348292 33794
rect 348240 33730 348292 33736
rect 347792 16546 348096 16574
rect 346768 15904 346820 15910
rect 346768 15846 346820 15852
rect 346412 6886 346992 6914
rect 346964 480 346992 6886
rect 348068 480 348096 16546
rect 349172 3346 349200 70994
rect 349264 58682 349292 84166
rect 349252 58676 349304 58682
rect 349252 58618 349304 58624
rect 349252 46300 349304 46306
rect 349252 46242 349304 46248
rect 349264 3466 349292 46242
rect 349448 26926 349476 96834
rect 349632 84194 349660 100028
rect 349712 96960 349764 96966
rect 349712 96902 349764 96908
rect 349540 84166 349660 84194
rect 349540 83502 349568 84166
rect 349528 83496 349580 83502
rect 349528 83438 349580 83444
rect 349724 54534 349752 96902
rect 349908 84194 349936 100028
rect 350092 96898 350120 100028
rect 350184 100014 350382 100042
rect 350184 96966 350212 100014
rect 350172 96960 350224 96966
rect 350172 96902 350224 96908
rect 350644 96898 350672 100028
rect 350828 97170 350856 100028
rect 350816 97164 350868 97170
rect 350816 97106 350868 97112
rect 350908 96960 350960 96966
rect 350908 96902 350960 96908
rect 350080 96892 350132 96898
rect 350080 96834 350132 96840
rect 350632 96892 350684 96898
rect 350632 96834 350684 96840
rect 349816 84166 349936 84194
rect 349816 71058 349844 84166
rect 349804 71052 349856 71058
rect 349804 70994 349856 71000
rect 349712 54528 349764 54534
rect 349712 54470 349764 54476
rect 349436 26920 349488 26926
rect 349436 26862 349488 26868
rect 350920 3466 350948 96902
rect 351104 93158 351132 100028
rect 351196 100014 351394 100042
rect 351196 96966 351224 100014
rect 351184 96960 351236 96966
rect 351184 96902 351236 96908
rect 351092 93152 351144 93158
rect 351092 93094 351144 93100
rect 351564 84194 351592 100028
rect 351196 84166 351592 84194
rect 351656 100014 351854 100042
rect 351196 3602 351224 84166
rect 351656 16574 351684 100014
rect 352564 97844 352616 97850
rect 352564 97786 352616 97792
rect 351920 93424 351972 93430
rect 351920 93366 351972 93372
rect 351656 16546 351776 16574
rect 351644 6248 351696 6254
rect 351644 6190 351696 6196
rect 351184 3596 351236 3602
rect 351184 3538 351236 3544
rect 349252 3460 349304 3466
rect 349252 3402 349304 3408
rect 350448 3460 350500 3466
rect 350448 3402 350500 3408
rect 350908 3460 350960 3466
rect 350908 3402 350960 3408
rect 349172 3318 349292 3346
rect 349264 480 349292 3318
rect 350460 480 350488 3402
rect 351656 480 351684 6190
rect 351748 3369 351776 16546
rect 351932 6914 351960 93366
rect 352576 11762 352604 97786
rect 352748 97028 352800 97034
rect 352748 96970 352800 96976
rect 352656 96892 352708 96898
rect 352656 96834 352708 96840
rect 352668 69698 352696 96834
rect 352760 73846 352788 96970
rect 352748 73840 352800 73846
rect 352748 73782 352800 73788
rect 352656 69692 352708 69698
rect 352656 69634 352708 69640
rect 353300 32496 353352 32502
rect 353300 32438 353352 32444
rect 353312 16574 353340 32438
rect 353312 16546 353616 16574
rect 352564 11756 352616 11762
rect 352564 11698 352616 11704
rect 351932 6886 352880 6914
rect 351734 3360 351790 3369
rect 351734 3295 351790 3304
rect 352852 480 352880 6886
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 353956 6866 353984 101759
rect 354048 20670 354076 105295
rect 354140 33114 354168 108831
rect 354232 46918 354260 112367
rect 354324 60722 354352 115903
rect 354416 73166 354444 119439
rect 354508 86970 354536 122975
rect 354600 100706 354628 126511
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 354588 100700 354640 100706
rect 354588 100642 354640 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 364984 97776 365036 97782
rect 364984 97718 365036 97724
rect 363604 97708 363656 97714
rect 363604 97650 363656 97656
rect 355324 97640 355376 97646
rect 355324 97582 355376 97588
rect 354496 86964 354548 86970
rect 354496 86906 354548 86912
rect 354404 73160 354456 73166
rect 354404 73102 354456 73108
rect 354312 60716 354364 60722
rect 354312 60658 354364 60664
rect 354220 46912 354272 46918
rect 354220 46854 354272 46860
rect 354128 33108 354180 33114
rect 354128 33050 354180 33056
rect 354680 31204 354732 31210
rect 354680 31146 354732 31152
rect 354036 20664 354088 20670
rect 354036 20606 354088 20612
rect 354692 16574 354720 31146
rect 354692 16546 355272 16574
rect 353944 6860 353996 6866
rect 353944 6802 353996 6808
rect 355244 480 355272 16546
rect 355336 9042 355364 97582
rect 360844 97572 360896 97578
rect 360844 97514 360896 97520
rect 355508 97504 355560 97510
rect 355508 97446 355560 97452
rect 355416 97164 355468 97170
rect 355416 97106 355468 97112
rect 355428 17270 355456 97106
rect 355520 83638 355548 97446
rect 356704 97436 356756 97442
rect 356704 97378 356756 97384
rect 356060 94784 356112 94790
rect 356060 94726 356112 94732
rect 355508 83632 355560 83638
rect 355508 83574 355560 83580
rect 355416 17264 355468 17270
rect 355416 17206 355468 17212
rect 356072 16574 356100 94726
rect 356072 16546 356376 16574
rect 355324 9036 355376 9042
rect 355324 8978 355376 8984
rect 356348 480 356376 16546
rect 356716 4894 356744 97378
rect 359464 97368 359516 97374
rect 359464 97310 359516 97316
rect 358820 91996 358872 92002
rect 358820 91938 358872 91944
rect 357440 74044 357492 74050
rect 357440 73986 357492 73992
rect 356704 4888 356756 4894
rect 356704 4830 356756 4836
rect 357452 3074 357480 73986
rect 357532 14476 357584 14482
rect 357532 14418 357584 14424
rect 357544 3194 357572 14418
rect 358832 6914 358860 91938
rect 359476 7682 359504 97310
rect 360200 72616 360252 72622
rect 360200 72558 360252 72564
rect 359464 7676 359516 7682
rect 359464 7618 359516 7624
rect 360212 6914 360240 72558
rect 360856 10402 360884 97514
rect 362960 90568 363012 90574
rect 362960 90510 363012 90516
rect 361580 61532 361632 61538
rect 361580 61474 361632 61480
rect 361592 16574 361620 61474
rect 362972 16574 363000 90510
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 360844 10396 360896 10402
rect 360844 10338 360896 10344
rect 358832 6886 359504 6914
rect 360212 6886 361160 6914
rect 357532 3188 357584 3194
rect 357532 3130 357584 3136
rect 358728 3188 358780 3194
rect 358728 3130 358780 3136
rect 357452 3046 357572 3074
rect 357544 480 357572 3046
rect 358740 480 358768 3130
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 6886
rect 361132 480 361160 6886
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 363616 13122 363644 97650
rect 364340 94716 364392 94722
rect 364340 94658 364392 94664
rect 364352 16574 364380 94658
rect 364352 16546 364656 16574
rect 363604 13116 363656 13122
rect 363604 13058 363656 13064
rect 364628 480 364656 16546
rect 364996 14482 365024 97718
rect 485044 97300 485096 97306
rect 485044 97242 485096 97248
rect 367100 96212 367152 96218
rect 367100 96154 367152 96160
rect 365720 86420 365772 86426
rect 365720 86362 365772 86368
rect 364984 14476 365036 14482
rect 364984 14418 365036 14424
rect 365732 1562 365760 86362
rect 365812 20052 365864 20058
rect 365812 19994 365864 20000
rect 365720 1556 365772 1562
rect 365720 1498 365772 1504
rect 365824 480 365852 19994
rect 367112 16574 367140 96154
rect 374000 96144 374052 96150
rect 374000 96086 374052 96092
rect 369860 89208 369912 89214
rect 369860 89150 369912 89156
rect 368480 85060 368532 85066
rect 368480 85002 368532 85008
rect 368492 16574 368520 85002
rect 369872 16574 369900 89150
rect 371240 80912 371292 80918
rect 371240 80854 371292 80860
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 367008 1556 367060 1562
rect 367008 1498 367060 1504
rect 367020 480 367048 1498
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 80854
rect 372620 62960 372672 62966
rect 372620 62902 372672 62908
rect 372632 16574 372660 62902
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3074 374040 96086
rect 431960 96076 432012 96082
rect 431960 96018 432012 96024
rect 386420 94648 386472 94654
rect 386420 94590 386472 94596
rect 376760 87848 376812 87854
rect 376760 87790 376812 87796
rect 374092 69828 374144 69834
rect 374092 69770 374144 69776
rect 374104 3194 374132 69770
rect 376772 16574 376800 87790
rect 383660 84992 383712 84998
rect 383660 84934 383712 84940
rect 380900 83700 380952 83706
rect 380900 83642 380952 83648
rect 378140 73976 378192 73982
rect 378140 73918 378192 73924
rect 378152 16574 378180 73918
rect 380912 16574 380940 83642
rect 382280 71188 382332 71194
rect 382280 71130 382332 71136
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 376024 13252 376076 13258
rect 376024 13194 376076 13200
rect 374092 3188 374144 3194
rect 374092 3130 374144 3136
rect 375288 3188 375340 3194
rect 375288 3130 375340 3136
rect 374012 3046 374132 3074
rect 374104 480 374132 3046
rect 375300 480 375328 3130
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 13194
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379520 11824 379572 11830
rect 379520 11766 379572 11772
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 11766
rect 381188 480 381216 16546
rect 382292 3074 382320 71130
rect 382372 26988 382424 26994
rect 382372 26930 382424 26936
rect 382384 3194 382412 26930
rect 383672 16574 383700 84934
rect 385040 72548 385092 72554
rect 385040 72490 385092 72496
rect 385052 16574 385080 72490
rect 386432 16574 386460 94590
rect 387800 93356 387852 93362
rect 387800 93298 387852 93304
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 382372 3188 382424 3194
rect 382372 3130 382424 3136
rect 383568 3188 383620 3194
rect 383568 3130 383620 3136
rect 382292 3046 382412 3074
rect 382384 480 382412 3046
rect 383580 480 383608 3130
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 93298
rect 390560 91928 390612 91934
rect 390560 91870 390612 91876
rect 389180 82272 389232 82278
rect 389180 82214 389232 82220
rect 389192 16574 389220 82214
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 1562 390600 91870
rect 394700 90500 394752 90506
rect 394700 90442 394752 90448
rect 391940 79484 391992 79490
rect 391940 79426 391992 79432
rect 390652 75336 390704 75342
rect 390652 75278 390704 75284
rect 390560 1556 390612 1562
rect 390560 1498 390612 1504
rect 390664 480 390692 75278
rect 391952 16574 391980 79426
rect 393320 17332 393372 17338
rect 393320 17274 393372 17280
rect 393332 16574 393360 17274
rect 394712 16574 394740 90442
rect 423680 89140 423732 89146
rect 423680 89082 423732 89088
rect 408500 86352 408552 86358
rect 408500 86294 408552 86300
rect 398840 80844 398892 80850
rect 398840 80786 398892 80792
rect 396080 60104 396132 60110
rect 396080 60046 396132 60052
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 391848 1556 391900 1562
rect 391848 1498 391900 1504
rect 391860 480 391888 1498
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 60046
rect 397736 6180 397788 6186
rect 397736 6122 397788 6128
rect 397748 480 397776 6122
rect 398852 3074 398880 80786
rect 401600 68468 401652 68474
rect 401600 68410 401652 68416
rect 400220 32428 400272 32434
rect 400220 32370 400272 32376
rect 398932 25628 398984 25634
rect 398932 25570 398984 25576
rect 398944 3194 398972 25570
rect 400232 16574 400260 32370
rect 401612 16574 401640 68410
rect 405740 67040 405792 67046
rect 405740 66982 405792 66988
rect 402980 57384 403032 57390
rect 402980 57326 403032 57332
rect 402992 16574 403020 57326
rect 404360 29708 404412 29714
rect 404360 29650 404412 29656
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 398932 3188 398984 3194
rect 398932 3130 398984 3136
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 398852 3046 398972 3074
rect 398944 480 398972 3046
rect 400140 480 400168 3130
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 29650
rect 405752 16574 405780 66982
rect 407120 64320 407172 64326
rect 407120 64262 407172 64268
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3194 407160 64262
rect 407212 24200 407264 24206
rect 407212 24142 407264 24148
rect 407120 3188 407172 3194
rect 407120 3130 407172 3136
rect 407224 480 407252 24142
rect 408512 16574 408540 86294
rect 409880 86284 409932 86290
rect 409880 86226 409932 86232
rect 409892 16574 409920 86226
rect 412640 82204 412692 82210
rect 412640 82146 412692 82152
rect 411260 28348 411312 28354
rect 411260 28290 411312 28296
rect 411272 16574 411300 28290
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 408420 480 408448 3130
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 82146
rect 415400 79416 415452 79422
rect 415400 79358 415452 79364
rect 414020 78124 414072 78130
rect 414020 78066 414072 78072
rect 414032 16574 414060 78066
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3194 415440 79358
rect 419540 65680 419592 65686
rect 419540 65622 419592 65628
rect 416780 56024 416832 56030
rect 416780 55966 416832 55972
rect 416792 16574 416820 55966
rect 418160 31136 418212 31142
rect 418160 31078 418212 31084
rect 418172 16574 418200 31078
rect 419552 16574 419580 65622
rect 422300 60036 422352 60042
rect 422300 59978 422352 59984
rect 420920 22840 420972 22846
rect 420920 22782 420972 22788
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 415492 14544 415544 14550
rect 415492 14486 415544 14492
rect 415400 3188 415452 3194
rect 415400 3130 415452 3136
rect 415504 480 415532 14486
rect 416688 3188 416740 3194
rect 416688 3130 416740 3136
rect 416700 480 416728 3130
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 22782
rect 422312 16574 422340 59978
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 3074 423720 89082
rect 430580 78056 430632 78062
rect 430580 77998 430632 78004
rect 426440 64252 426492 64258
rect 426440 64194 426492 64200
rect 423772 21480 423824 21486
rect 423772 21422 423824 21428
rect 423784 3194 423812 21422
rect 425060 19984 425112 19990
rect 425060 19926 425112 19932
rect 425072 16574 425100 19926
rect 426452 16574 426480 64194
rect 427820 54664 427872 54670
rect 427820 54606 427872 54612
rect 427832 16574 427860 54606
rect 430592 16574 430620 77998
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 423772 3188 423824 3194
rect 423772 3130 423824 3136
rect 424968 3188 425020 3194
rect 424968 3130 425020 3136
rect 423692 3046 423812 3074
rect 423784 480 423812 3046
rect 424980 480 425008 3130
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429200 13184 429252 13190
rect 429200 13126 429252 13132
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 13126
rect 430868 480 430896 16546
rect 431972 3194 432000 96018
rect 458180 93288 458232 93294
rect 458180 93230 458232 93236
rect 452660 89072 452712 89078
rect 452660 89014 452712 89020
rect 440332 87780 440384 87786
rect 440332 87722 440384 87728
rect 434720 69760 434772 69766
rect 434720 69702 434772 69708
rect 433340 62892 433392 62898
rect 433340 62834 433392 62840
rect 432052 18692 432104 18698
rect 432052 18634 432104 18640
rect 431960 3188 432012 3194
rect 431960 3130 432012 3136
rect 432064 480 432092 18634
rect 433352 16574 433380 62834
rect 434732 16574 434760 69702
rect 437480 61464 437532 61470
rect 437480 61406 437532 61412
rect 436100 58812 436152 58818
rect 436100 58754 436152 58760
rect 436112 16574 436140 58754
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433248 3188 433300 3194
rect 433248 3130 433300 3136
rect 433260 480 433288 3130
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 61406
rect 438860 51808 438912 51814
rect 438860 51750 438912 51756
rect 438872 16574 438900 51750
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440344 3262 440372 87722
rect 448520 76696 448572 76702
rect 448520 76638 448572 76644
rect 441620 73908 441672 73914
rect 441620 73850 441672 73856
rect 441632 16574 441660 73850
rect 444380 58744 444432 58750
rect 444380 58686 444432 58692
rect 444392 16574 444420 58686
rect 445760 50448 445812 50454
rect 445760 50390 445812 50396
rect 441632 16546 442672 16574
rect 444392 16546 445064 16574
rect 440240 3256 440292 3262
rect 440240 3198 440292 3204
rect 440332 3256 440384 3262
rect 440332 3198 440384 3204
rect 441528 3256 441580 3262
rect 441528 3198 441580 3204
rect 440252 1714 440280 3198
rect 440252 1686 440372 1714
rect 440344 480 440372 1686
rect 441540 480 441568 3198
rect 442644 480 442672 16546
rect 443828 3324 443880 3330
rect 443828 3266 443880 3272
rect 443840 480 443868 3266
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 50390
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 447428 480 447456 3334
rect 448532 3210 448560 76638
rect 451280 57316 451332 57322
rect 451280 57258 451332 57264
rect 448612 53168 448664 53174
rect 448612 53110 448664 53116
rect 448624 3398 448652 53110
rect 451292 16574 451320 57258
rect 452672 16574 452700 89014
rect 455420 83564 455472 83570
rect 455420 83506 455472 83512
rect 455432 16574 455460 83506
rect 456892 71120 456944 71126
rect 456892 71062 456944 71068
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 455432 16546 455736 16574
rect 450912 4140 450964 4146
rect 450912 4082 450964 4088
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 4082
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 454500 4072 454552 4078
rect 454500 4014 454552 4020
rect 454512 480 454540 4014
rect 455708 480 455736 16546
rect 456904 480 456932 71062
rect 458192 16574 458220 93230
rect 477500 87712 477552 87718
rect 477500 87654 477552 87660
rect 459560 80776 459612 80782
rect 459560 80718 459612 80724
rect 459572 16574 459600 80718
rect 470600 72480 470652 72486
rect 470600 72422 470652 72428
rect 462320 55956 462372 55962
rect 462320 55898 462372 55904
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 458088 4004 458140 4010
rect 458088 3946 458140 3952
rect 458100 480 458128 3946
rect 459204 480 459232 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 461596 480 461624 3878
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 55898
rect 465172 54596 465224 54602
rect 465172 54538 465224 54544
rect 463700 25560 463752 25566
rect 463700 25502 463752 25508
rect 463712 16574 463740 25502
rect 465184 16574 465212 54538
rect 469220 53100 469272 53106
rect 469220 53042 469272 53048
rect 466460 24132 466512 24138
rect 466460 24074 466512 24080
rect 466472 16574 466500 24074
rect 469232 16574 469260 53042
rect 463712 16546 464016 16574
rect 465184 16546 465856 16574
rect 466472 16546 467512 16574
rect 469232 16546 469904 16574
rect 463988 480 464016 16546
rect 465172 3868 465224 3874
rect 465172 3810 465224 3816
rect 465184 480 465212 3810
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 468668 3800 468720 3806
rect 468668 3742 468720 3748
rect 468680 480 468708 3742
rect 469876 480 469904 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 72422
rect 476120 68400 476172 68406
rect 476120 68342 476172 68348
rect 473360 51740 473412 51746
rect 473360 51682 473412 51688
rect 473372 6914 473400 51682
rect 473452 22772 473504 22778
rect 473452 22714 473504 22720
rect 473464 16574 473492 22714
rect 476132 16574 476160 68342
rect 477512 16574 477540 87654
rect 480260 83632 480312 83638
rect 480260 83574 480312 83580
rect 480272 16574 480300 83574
rect 481640 75268 481692 75274
rect 481640 75210 481692 75216
rect 473464 16546 474136 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 473372 6886 473492 6914
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473464 480 473492 6886
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475764 480 475792 3606
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481652 6914 481680 75210
rect 484400 50380 484452 50386
rect 484400 50322 484452 50328
rect 481732 49088 481784 49094
rect 481732 49030 481784 49036
rect 481744 16574 481772 49030
rect 484412 16574 484440 50322
rect 481744 16546 482416 16574
rect 484412 16546 484808 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484032 4888 484084 4894
rect 484032 4830 484084 4836
rect 484044 480 484072 4830
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 485056 4214 485084 97242
rect 489920 96008 489972 96014
rect 489920 95950 489972 95956
rect 485780 76628 485832 76634
rect 485780 76570 485832 76576
rect 485792 16574 485820 76570
rect 488540 66972 488592 66978
rect 488540 66914 488592 66920
rect 488552 16574 488580 66914
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 485044 4208 485096 4214
rect 485044 4150 485096 4156
rect 486436 480 486464 16546
rect 487620 4208 487672 4214
rect 487620 4150 487672 4156
rect 487632 480 487660 4150
rect 488828 480 488856 16546
rect 489932 3534 489960 95950
rect 543740 95940 543792 95946
rect 543740 95882 543792 95888
rect 494060 94580 494112 94586
rect 494060 94522 494112 94528
rect 491300 49020 491352 49026
rect 491300 48962 491352 48968
rect 490012 21412 490064 21418
rect 490012 21354 490064 21360
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 21354
rect 491312 16574 491340 48962
rect 492680 18624 492732 18630
rect 492680 18566 492732 18572
rect 492692 16574 492720 18566
rect 494072 16574 494100 94522
rect 498200 93220 498252 93226
rect 498200 93162 498252 93168
rect 495440 65612 495492 65618
rect 495440 65554 495492 65560
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 65554
rect 497096 4820 497148 4826
rect 497096 4762 497148 4768
rect 497108 480 497136 4762
rect 498212 480 498240 93162
rect 507860 91860 507912 91866
rect 507860 91802 507912 91808
rect 503720 68332 503772 68338
rect 503720 68274 503772 68280
rect 498292 47660 498344 47666
rect 498292 47602 498344 47608
rect 498304 16574 498332 47602
rect 499580 46232 499632 46238
rect 499580 46174 499632 46180
rect 499592 16574 499620 46174
rect 502340 44940 502392 44946
rect 502340 44882 502392 44888
rect 502352 16574 502380 44882
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 501788 7676 501840 7682
rect 501788 7618 501840 7624
rect 501800 480 501828 7618
rect 502996 480 503024 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 68274
rect 506480 43512 506532 43518
rect 506480 43454 506532 43460
rect 505376 9036 505428 9042
rect 505376 8978 505428 8984
rect 505388 480 505416 8978
rect 506492 480 506520 43454
rect 507872 16574 507900 91802
rect 512000 90432 512052 90438
rect 512000 90374 512052 90380
rect 510620 47592 510672 47598
rect 510620 47534 510672 47540
rect 509240 42152 509292 42158
rect 509240 42094 509292 42100
rect 509252 16574 509280 42094
rect 510632 16574 510660 47534
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 507676 7608 507728 7614
rect 507676 7550 507728 7556
rect 507688 480 507716 7550
rect 508884 480 508912 16546
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 90374
rect 518900 89004 518952 89010
rect 518900 88946 518952 88952
rect 517520 57248 517572 57254
rect 517520 57190 517572 57196
rect 513380 40792 513432 40798
rect 513380 40734 513432 40740
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 40734
rect 516140 39432 516192 39438
rect 516140 39374 516192 39380
rect 516152 16574 516180 39374
rect 517532 16574 517560 57190
rect 518912 16574 518940 88946
rect 523040 87644 523092 87650
rect 523040 87586 523092 87592
rect 521660 44872 521712 44878
rect 521660 44814 521712 44820
rect 520280 38004 520332 38010
rect 520280 37946 520332 37952
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515496 10396 515548 10402
rect 515496 10338 515548 10344
rect 514760 8968 514812 8974
rect 514760 8910 514812 8916
rect 514772 480 514800 8910
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 10338
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 37946
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 44814
rect 523052 480 523080 87586
rect 525800 84924 525852 84930
rect 525800 84866 525852 84872
rect 524420 43444 524472 43450
rect 524420 43386 524472 43392
rect 524432 16574 524460 43386
rect 525812 16574 525840 84866
rect 529940 82136 529992 82142
rect 529940 82078 529992 82084
rect 528560 42084 528612 42090
rect 528560 42026 528612 42032
rect 527180 36644 527232 36650
rect 527180 36586 527232 36592
rect 527192 16574 527220 36586
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523776 15972 523828 15978
rect 523776 15914 523828 15920
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 15914
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 42026
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 82078
rect 536840 80708 536892 80714
rect 536840 80650 536892 80656
rect 535460 66904 535512 66910
rect 535460 66846 535512 66852
rect 531320 64184 531372 64190
rect 531320 64126 531372 64132
rect 531332 480 531360 64126
rect 534080 35284 534132 35290
rect 534080 35226 534132 35232
rect 534092 16574 534120 35226
rect 535472 16574 535500 66846
rect 536852 16574 536880 80650
rect 539600 79348 539652 79354
rect 539600 79290 539652 79296
rect 538220 33856 538272 33862
rect 538220 33798 538272 33804
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 533712 11756 533764 11762
rect 533712 11698 533764 11704
rect 532056 10328 532108 10334
rect 532056 10270 532108 10276
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 10270
rect 533724 480 533752 11698
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 33798
rect 539612 3534 539640 79290
rect 542360 55888 542412 55894
rect 542360 55830 542412 55836
rect 539692 40724 539744 40730
rect 539692 40666 539744 40672
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 40666
rect 540980 31068 541032 31074
rect 540980 31010 541032 31016
rect 540992 16574 541020 31010
rect 542372 16574 542400 55830
rect 543752 16574 543780 95882
rect 557540 94512 557592 94518
rect 557540 94454 557592 94460
rect 545120 91792 545172 91798
rect 545120 91734 545172 91740
rect 545132 16574 545160 91734
rect 547880 77988 547932 77994
rect 547880 77930 547932 77936
rect 546500 39364 546552 39370
rect 546500 39306 546552 39312
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 39306
rect 547892 480 547920 77930
rect 554780 76560 554832 76566
rect 554780 76502 554832 76508
rect 552020 62824 552072 62830
rect 552020 62766 552072 62772
rect 549260 37936 549312 37942
rect 549260 37878 549312 37884
rect 547972 29640 548024 29646
rect 547972 29582 548024 29588
rect 547984 16574 548012 29582
rect 549272 16574 549300 37878
rect 552032 16574 552060 62766
rect 553400 36576 553452 36582
rect 553400 36518 553452 36524
rect 553412 16574 553440 36518
rect 547984 16546 548656 16574
rect 549272 16546 550312 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 551008 13116 551060 13122
rect 551008 13058 551060 13064
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 13058
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 76502
rect 556160 61396 556212 61402
rect 556160 61338 556212 61344
rect 556172 480 556200 61338
rect 556252 35216 556304 35222
rect 556252 35158 556304 35164
rect 556264 16574 556292 35158
rect 557552 16574 557580 94454
rect 578240 93152 578292 93158
rect 578240 93094 578292 93100
rect 563060 90364 563112 90370
rect 563060 90306 563112 90312
rect 561680 75200 561732 75206
rect 561680 75142 561732 75148
rect 558920 28280 558972 28286
rect 558920 28222 558972 28228
rect 558932 16574 558960 28222
rect 561692 16574 561720 75142
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 560392 15904 560444 15910
rect 560392 15846 560444 15852
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 15846
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 90306
rect 565820 84856 565872 84862
rect 565820 84798 565872 84804
rect 564532 73840 564584 73846
rect 564532 73782 564584 73788
rect 563704 65544 563756 65550
rect 563704 65486 563756 65492
rect 563716 3534 563744 65486
rect 564544 16574 564572 73782
rect 565832 16574 565860 84798
rect 571340 83496 571392 83502
rect 571340 83438 571392 83444
rect 569960 58676 570012 58682
rect 569960 58618 570012 58624
rect 567200 33788 567252 33794
rect 567200 33730 567252 33736
rect 567212 16574 567240 33730
rect 569972 16574 570000 58618
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 563704 3528 563756 3534
rect 563704 3470 563756 3476
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564452 480 564480 3470
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 568672 14476 568724 14482
rect 568672 14418 568724 14424
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 14418
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 83438
rect 571984 71052 572036 71058
rect 571984 70994 572036 71000
rect 571996 3534 572024 70994
rect 575480 69692 575532 69698
rect 575480 69634 575532 69640
rect 574100 54528 574152 54534
rect 574100 54470 574152 54476
rect 572812 26920 572864 26926
rect 572812 26862 572864 26868
rect 572824 16574 572852 26862
rect 574112 16574 574140 54470
rect 575492 16574 575520 69634
rect 576860 17264 576912 17270
rect 576860 17206 576912 17212
rect 576872 16574 576900 17206
rect 578252 16574 578280 93094
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 572824 16546 573496 16574
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 572732 480 572760 3470
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3422 671200 3478 671256
rect 3330 632068 3332 632088
rect 3332 632068 3384 632088
rect 3384 632068 3386 632088
rect 3330 632032 3386 632068
rect 3330 619112 3386 619168
rect 3330 606056 3386 606112
rect 3146 579944 3202 580000
rect 2962 527856 3018 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3238 501744 3294 501800
rect 3330 475632 3386 475688
rect 2962 423544 3018 423600
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3146 319232 3202 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 3238 267144 3294 267200
rect 3514 658144 3570 658200
rect 3330 254088 3386 254144
rect 3606 566888 3662 566944
rect 3422 241032 3478 241088
rect 3698 553832 3754 553888
rect 3790 462576 3846 462632
rect 3514 214920 3570 214976
rect 3882 449520 3938 449576
rect 3974 358400 4030 358456
rect 3606 201864 3662 201920
rect 3698 188808 3754 188864
rect 3422 149776 3478 149832
rect 4066 345344 4122 345400
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 229098 258032 229154 258088
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 353942 254496 353998 254552
rect 229466 254224 229522 254280
rect 353298 250960 353354 251016
rect 230386 250416 230442 250472
rect 353298 247424 353354 247480
rect 229834 246608 229890 246664
rect 353298 243888 353354 243944
rect 229650 242836 229652 242856
rect 229652 242836 229704 242856
rect 229704 242836 229706 242856
rect 229650 242800 229706 242836
rect 353298 240352 353354 240408
rect 230386 238992 230442 239048
rect 353298 236816 353354 236872
rect 229834 235184 229890 235240
rect 353298 233180 353300 233200
rect 353300 233180 353352 233200
rect 353352 233180 353354 233200
rect 353298 233144 353354 233180
rect 230386 231376 230442 231432
rect 353298 229608 353354 229664
rect 230386 227568 230442 227624
rect 353298 226072 353354 226128
rect 230386 223760 230442 223816
rect 353298 222536 353354 222592
rect 230386 219952 230442 220008
rect 353298 219000 353354 219056
rect 230386 216144 230442 216200
rect 353298 215464 353354 215520
rect 230386 212336 230442 212392
rect 353298 211928 353354 211984
rect 230018 208528 230074 208584
rect 353298 208392 353354 208448
rect 230386 204720 230442 204776
rect 353298 204720 353354 204776
rect 353298 201184 353354 201240
rect 229650 200912 229706 200968
rect 353298 197648 353354 197704
rect 230386 197104 230442 197160
rect 353298 194112 353354 194168
rect 229650 193296 229706 193352
rect 230386 189488 230442 189544
rect 353298 187040 353354 187096
rect 230386 185680 230442 185736
rect 353298 183524 353354 183560
rect 353298 183504 353300 183524
rect 353300 183504 353352 183524
rect 353352 183504 353354 183524
rect 230386 181872 230442 181928
rect 353298 179832 353354 179888
rect 229650 178064 229706 178120
rect 353298 176296 353354 176352
rect 230386 174256 230442 174312
rect 353298 172760 353354 172816
rect 230386 170448 230442 170504
rect 230386 166640 230442 166696
rect 353298 165688 353354 165744
rect 3790 162832 3846 162888
rect 229650 162832 229706 162888
rect 353298 162152 353354 162208
rect 229466 159024 229522 159080
rect 354310 258168 354366 258224
rect 354034 190576 354090 190632
rect 353942 158616 353998 158672
rect 230386 155216 230442 155272
rect 353298 155080 353354 155136
rect 230386 151408 230442 151464
rect 353298 151408 353354 151464
rect 229650 147620 229706 147656
rect 229650 147600 229652 147620
rect 229652 147600 229704 147620
rect 229704 147600 229706 147620
rect 353298 144336 353354 144392
rect 230386 143792 230442 143848
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 365064 580226 365120
rect 579986 325216 580042 325272
rect 579802 312024 579858 312080
rect 580170 298696 580226 298752
rect 354126 169224 354182 169280
rect 580354 590960 580410 591016
rect 580170 258848 580226 258904
rect 580170 245520 580226 245576
rect 580446 577632 580502 577688
rect 580538 484608 580594 484664
rect 580262 232328 580318 232384
rect 580170 219000 580226 219056
rect 580170 179152 580226 179208
rect 580630 471416 580686 471472
rect 580722 378392 580778 378448
rect 580354 205672 580410 205728
rect 580814 351872 580870 351928
rect 580446 192480 580502 192536
rect 580170 152632 580226 152688
rect 580906 272176 580962 272232
rect 580538 165824 580594 165880
rect 354034 147872 354090 147928
rect 353942 140800 353998 140856
rect 230386 139984 230442 140040
rect 580170 139304 580226 139360
rect 353298 137264 353354 137320
rect 3422 136720 3478 136776
rect 229834 136176 229890 136232
rect 354310 133728 354366 133784
rect 229742 132368 229798 132424
rect 3146 110608 3202 110664
rect 3330 84632 3386 84688
rect 3330 71576 3386 71632
rect 353942 130192 353998 130248
rect 230386 128560 230442 128616
rect 230110 124752 230166 124808
rect 230018 120944 230074 121000
rect 229926 113328 229982 113384
rect 229834 109520 229890 109576
rect 229742 101904 229798 101960
rect 3606 97552 3662 97608
rect 3514 58520 3570 58576
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 6458 3304 6514 3360
rect 230202 117136 230258 117192
rect 354586 126520 354642 126576
rect 354494 122984 354550 123040
rect 354402 119448 354458 119504
rect 354310 115912 354366 115968
rect 354218 112376 354274 112432
rect 354126 108840 354182 108896
rect 230386 105712 230442 105768
rect 354034 105304 354090 105360
rect 353942 101768 353998 101824
rect 233330 3304 233386 3360
rect 351734 3304 351790 3360
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 580441 577690 580507 577693
rect 583520 577690 584960 577780
rect 580441 577688 584960 577690
rect 580441 577632 580446 577688
rect 580502 577632 584960 577688
rect 580441 577630 584960 577632
rect 580441 577627 580507 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580625 471474 580691 471477
rect 583520 471474 584960 471564
rect 580625 471472 584960 471474
rect 580625 471416 580630 471472
rect 580686 471416 584960 471472
rect 580625 471414 584960 471416
rect 580625 471411 580691 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3785 462634 3851 462637
rect -960 462632 3851 462634
rect -960 462576 3790 462632
rect 3846 462576 3851 462632
rect -960 462574 3851 462576
rect -960 462484 480 462574
rect 3785 462571 3851 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3877 449578 3943 449581
rect -960 449576 3943 449578
rect -960 449520 3882 449576
rect 3938 449520 3943 449576
rect -960 449518 3943 449520
rect -960 449428 480 449518
rect 3877 449515 3943 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2957 423602 3023 423605
rect -960 423600 3023 423602
rect -960 423544 2962 423600
rect 3018 423544 3023 423600
rect -960 423542 3023 423544
rect -960 423452 480 423542
rect 2957 423539 3023 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580717 378450 580783 378453
rect 583520 378450 584960 378540
rect 580717 378448 584960 378450
rect 580717 378392 580722 378448
rect 580778 378392 584960 378448
rect 580717 378390 584960 378392
rect 580717 378387 580783 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3969 358458 4035 358461
rect -960 358456 4035 358458
rect -960 358400 3974 358456
rect 4030 358400 4035 358456
rect -960 358398 4035 358400
rect -960 358308 480 358398
rect 3969 358395 4035 358398
rect 580809 351930 580875 351933
rect 583520 351930 584960 352020
rect 580809 351928 584960 351930
rect 580809 351872 580814 351928
rect 580870 351872 584960 351928
rect 580809 351870 584960 351872
rect 580809 351867 580875 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 4061 345402 4127 345405
rect -960 345400 4127 345402
rect -960 345344 4066 345400
rect 4122 345344 4127 345400
rect -960 345342 4127 345344
rect -960 345252 480 345342
rect 4061 345339 4127 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 579797 312082 579863 312085
rect 583520 312082 584960 312172
rect 579797 312080 584960 312082
rect 579797 312024 579802 312080
rect 579858 312024 584960 312080
rect 579797 312022 584960 312024
rect 579797 312019 579863 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580901 272234 580967 272237
rect 583520 272234 584960 272324
rect 580901 272232 584960 272234
rect 580901 272176 580906 272232
rect 580962 272176 584960 272232
rect 580901 272174 584960 272176
rect 580901 272171 580967 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 354305 258226 354371 258229
rect 354078 258224 354371 258226
rect 354078 258168 354310 258224
rect 354366 258168 354371 258224
rect 354078 258166 354371 258168
rect 229093 258090 229159 258093
rect 229093 258088 229202 258090
rect 229093 258032 229098 258088
rect 229154 258032 229202 258088
rect 229093 258027 229202 258032
rect 229142 257954 229202 258027
rect 231534 258030 232116 258090
rect 351900 258030 352482 258090
rect 231534 257954 231594 258030
rect 229142 257894 231594 257954
rect 352422 257954 352482 258030
rect 354078 257954 354138 258166
rect 354305 258163 354371 258166
rect 352422 257894 354138 257954
rect 353937 254554 354003 254557
rect 351900 254552 354003 254554
rect 351900 254496 353942 254552
rect 353998 254496 354003 254552
rect 351900 254494 354003 254496
rect 353937 254491 354003 254494
rect 229461 254282 229527 254285
rect 229461 254280 232116 254282
rect -960 254146 480 254236
rect 229461 254224 229466 254280
rect 229522 254224 232116 254280
rect 229461 254222 232116 254224
rect 229461 254219 229527 254222
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 353293 251018 353359 251021
rect 351900 251016 353359 251018
rect 351900 250960 353298 251016
rect 353354 250960 353359 251016
rect 351900 250958 353359 250960
rect 353293 250955 353359 250958
rect 230381 250474 230447 250477
rect 230381 250472 232116 250474
rect 230381 250416 230386 250472
rect 230442 250416 232116 250472
rect 230381 250414 232116 250416
rect 230381 250411 230447 250414
rect 353293 247482 353359 247485
rect 351900 247480 353359 247482
rect 351900 247424 353298 247480
rect 353354 247424 353359 247480
rect 351900 247422 353359 247424
rect 353293 247419 353359 247422
rect 229829 246666 229895 246669
rect 229829 246664 232116 246666
rect 229829 246608 229834 246664
rect 229890 246608 232116 246664
rect 229829 246606 232116 246608
rect 229829 246603 229895 246606
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 353293 243946 353359 243949
rect 351900 243944 353359 243946
rect 351900 243888 353298 243944
rect 353354 243888 353359 243944
rect 351900 243886 353359 243888
rect 353293 243883 353359 243886
rect 229645 242858 229711 242861
rect 229645 242856 232116 242858
rect 229645 242800 229650 242856
rect 229706 242800 232116 242856
rect 229645 242798 232116 242800
rect 229645 242795 229711 242798
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 353293 240410 353359 240413
rect 351900 240408 353359 240410
rect 351900 240352 353298 240408
rect 353354 240352 353359 240408
rect 351900 240350 353359 240352
rect 353293 240347 353359 240350
rect 230381 239050 230447 239053
rect 230381 239048 232116 239050
rect 230381 238992 230386 239048
rect 230442 238992 232116 239048
rect 230381 238990 232116 238992
rect 230381 238987 230447 238990
rect 353293 236874 353359 236877
rect 351900 236872 353359 236874
rect 351900 236816 353298 236872
rect 353354 236816 353359 236872
rect 351900 236814 353359 236816
rect 353293 236811 353359 236814
rect 229829 235242 229895 235245
rect 229829 235240 232116 235242
rect 229829 235184 229834 235240
rect 229890 235184 232116 235240
rect 229829 235182 232116 235184
rect 229829 235179 229895 235182
rect 353293 233202 353359 233205
rect 351900 233200 353359 233202
rect 351900 233144 353298 233200
rect 353354 233144 353359 233200
rect 351900 233142 353359 233144
rect 353293 233139 353359 233142
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect 230381 231434 230447 231437
rect 230381 231432 232116 231434
rect 230381 231376 230386 231432
rect 230442 231376 232116 231432
rect 230381 231374 232116 231376
rect 230381 231371 230447 231374
rect 353293 229666 353359 229669
rect 351900 229664 353359 229666
rect 351900 229608 353298 229664
rect 353354 229608 353359 229664
rect 351900 229606 353359 229608
rect 353293 229603 353359 229606
rect -960 227884 480 228124
rect 230381 227626 230447 227629
rect 230381 227624 232116 227626
rect 230381 227568 230386 227624
rect 230442 227568 232116 227624
rect 230381 227566 232116 227568
rect 230381 227563 230447 227566
rect 353293 226130 353359 226133
rect 351900 226128 353359 226130
rect 351900 226072 353298 226128
rect 353354 226072 353359 226128
rect 351900 226070 353359 226072
rect 353293 226067 353359 226070
rect 230381 223818 230447 223821
rect 230381 223816 232116 223818
rect 230381 223760 230386 223816
rect 230442 223760 232116 223816
rect 230381 223758 232116 223760
rect 230381 223755 230447 223758
rect 353293 222594 353359 222597
rect 351900 222592 353359 222594
rect 351900 222536 353298 222592
rect 353354 222536 353359 222592
rect 351900 222534 353359 222536
rect 353293 222531 353359 222534
rect 230381 220010 230447 220013
rect 230381 220008 232116 220010
rect 230381 219952 230386 220008
rect 230442 219952 232116 220008
rect 230381 219950 232116 219952
rect 230381 219947 230447 219950
rect 353293 219058 353359 219061
rect 351900 219056 353359 219058
rect 351900 219000 353298 219056
rect 353354 219000 353359 219056
rect 351900 218998 353359 219000
rect 353293 218995 353359 218998
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 230381 216202 230447 216205
rect 230381 216200 232116 216202
rect 230381 216144 230386 216200
rect 230442 216144 232116 216200
rect 230381 216142 232116 216144
rect 230381 216139 230447 216142
rect 353293 215522 353359 215525
rect 351900 215520 353359 215522
rect 351900 215464 353298 215520
rect 353354 215464 353359 215520
rect 351900 215462 353359 215464
rect 353293 215459 353359 215462
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 230381 212394 230447 212397
rect 230381 212392 232116 212394
rect 230381 212336 230386 212392
rect 230442 212336 232116 212392
rect 230381 212334 232116 212336
rect 230381 212331 230447 212334
rect 353293 211986 353359 211989
rect 351900 211984 353359 211986
rect 351900 211928 353298 211984
rect 353354 211928 353359 211984
rect 351900 211926 353359 211928
rect 353293 211923 353359 211926
rect 230013 208586 230079 208589
rect 230013 208584 232116 208586
rect 230013 208528 230018 208584
rect 230074 208528 232116 208584
rect 230013 208526 232116 208528
rect 230013 208523 230079 208526
rect 353293 208450 353359 208453
rect 351900 208448 353359 208450
rect 351900 208392 353298 208448
rect 353354 208392 353359 208448
rect 351900 208390 353359 208392
rect 353293 208387 353359 208390
rect 580349 205730 580415 205733
rect 583520 205730 584960 205820
rect 580349 205728 584960 205730
rect 580349 205672 580354 205728
rect 580410 205672 584960 205728
rect 580349 205670 584960 205672
rect 580349 205667 580415 205670
rect 583520 205580 584960 205670
rect 230381 204778 230447 204781
rect 353293 204778 353359 204781
rect 230381 204776 232116 204778
rect 230381 204720 230386 204776
rect 230442 204720 232116 204776
rect 230381 204718 232116 204720
rect 351900 204776 353359 204778
rect 351900 204720 353298 204776
rect 353354 204720 353359 204776
rect 351900 204718 353359 204720
rect 230381 204715 230447 204718
rect 353293 204715 353359 204718
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 353293 201242 353359 201245
rect 351900 201240 353359 201242
rect 351900 201184 353298 201240
rect 353354 201184 353359 201240
rect 351900 201182 353359 201184
rect 353293 201179 353359 201182
rect 229645 200970 229711 200973
rect 229645 200968 232116 200970
rect 229645 200912 229650 200968
rect 229706 200912 232116 200968
rect 229645 200910 232116 200912
rect 229645 200907 229711 200910
rect 353293 197706 353359 197709
rect 351900 197704 353359 197706
rect 351900 197648 353298 197704
rect 353354 197648 353359 197704
rect 351900 197646 353359 197648
rect 353293 197643 353359 197646
rect 230381 197162 230447 197165
rect 230381 197160 232116 197162
rect 230381 197104 230386 197160
rect 230442 197104 232116 197160
rect 230381 197102 232116 197104
rect 230381 197099 230447 197102
rect 353293 194170 353359 194173
rect 351900 194168 353359 194170
rect 351900 194112 353298 194168
rect 353354 194112 353359 194168
rect 351900 194110 353359 194112
rect 353293 194107 353359 194110
rect 229645 193354 229711 193357
rect 229645 193352 232116 193354
rect 229645 193296 229650 193352
rect 229706 193296 232116 193352
rect 229645 193294 232116 193296
rect 229645 193291 229711 193294
rect 580441 192538 580507 192541
rect 583520 192538 584960 192628
rect 580441 192536 584960 192538
rect 580441 192480 580446 192536
rect 580502 192480 584960 192536
rect 580441 192478 584960 192480
rect 580441 192475 580507 192478
rect 583520 192388 584960 192478
rect 354029 190634 354095 190637
rect 351900 190632 354095 190634
rect 351900 190576 354034 190632
rect 354090 190576 354095 190632
rect 351900 190574 354095 190576
rect 354029 190571 354095 190574
rect 230381 189546 230447 189549
rect 230381 189544 232116 189546
rect 230381 189488 230386 189544
rect 230442 189488 232116 189544
rect 230381 189486 232116 189488
rect 230381 189483 230447 189486
rect -960 188866 480 188956
rect 3693 188866 3759 188869
rect -960 188864 3759 188866
rect -960 188808 3698 188864
rect 3754 188808 3759 188864
rect -960 188806 3759 188808
rect -960 188716 480 188806
rect 3693 188803 3759 188806
rect 353293 187098 353359 187101
rect 351900 187096 353359 187098
rect 351900 187040 353298 187096
rect 353354 187040 353359 187096
rect 351900 187038 353359 187040
rect 353293 187035 353359 187038
rect 230381 185738 230447 185741
rect 230381 185736 232116 185738
rect 230381 185680 230386 185736
rect 230442 185680 232116 185736
rect 230381 185678 232116 185680
rect 230381 185675 230447 185678
rect 353293 183562 353359 183565
rect 351900 183560 353359 183562
rect 351900 183504 353298 183560
rect 353354 183504 353359 183560
rect 351900 183502 353359 183504
rect 353293 183499 353359 183502
rect 230381 181930 230447 181933
rect 230381 181928 232116 181930
rect 230381 181872 230386 181928
rect 230442 181872 232116 181928
rect 230381 181870 232116 181872
rect 230381 181867 230447 181870
rect 353293 179890 353359 179893
rect 351900 179888 353359 179890
rect 351900 179832 353298 179888
rect 353354 179832 353359 179888
rect 351900 179830 353359 179832
rect 353293 179827 353359 179830
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 229645 178122 229711 178125
rect 229645 178120 232116 178122
rect 229645 178064 229650 178120
rect 229706 178064 232116 178120
rect 229645 178062 232116 178064
rect 229645 178059 229711 178062
rect 353293 176354 353359 176357
rect 351900 176352 353359 176354
rect 351900 176296 353298 176352
rect 353354 176296 353359 176352
rect 351900 176294 353359 176296
rect 353293 176291 353359 176294
rect -960 175796 480 176036
rect 230381 174314 230447 174317
rect 230381 174312 232116 174314
rect 230381 174256 230386 174312
rect 230442 174256 232116 174312
rect 230381 174254 232116 174256
rect 230381 174251 230447 174254
rect 353293 172818 353359 172821
rect 351900 172816 353359 172818
rect 351900 172760 353298 172816
rect 353354 172760 353359 172816
rect 351900 172758 353359 172760
rect 353293 172755 353359 172758
rect 230381 170506 230447 170509
rect 230381 170504 232116 170506
rect 230381 170448 230386 170504
rect 230442 170448 232116 170504
rect 230381 170446 232116 170448
rect 230381 170443 230447 170446
rect 354121 169282 354187 169285
rect 351900 169280 354187 169282
rect 351900 169224 354126 169280
rect 354182 169224 354187 169280
rect 351900 169222 354187 169224
rect 354121 169219 354187 169222
rect 230381 166698 230447 166701
rect 230381 166696 232116 166698
rect 230381 166640 230386 166696
rect 230442 166640 232116 166696
rect 230381 166638 232116 166640
rect 230381 166635 230447 166638
rect 580533 165882 580599 165885
rect 583520 165882 584960 165972
rect 580533 165880 584960 165882
rect 580533 165824 580538 165880
rect 580594 165824 584960 165880
rect 580533 165822 584960 165824
rect 580533 165819 580599 165822
rect 353293 165746 353359 165749
rect 351900 165744 353359 165746
rect 351900 165688 353298 165744
rect 353354 165688 353359 165744
rect 583520 165732 584960 165822
rect 351900 165686 353359 165688
rect 353293 165683 353359 165686
rect -960 162890 480 162980
rect 3785 162890 3851 162893
rect -960 162888 3851 162890
rect -960 162832 3790 162888
rect 3846 162832 3851 162888
rect -960 162830 3851 162832
rect -960 162740 480 162830
rect 3785 162827 3851 162830
rect 229645 162890 229711 162893
rect 229645 162888 232116 162890
rect 229645 162832 229650 162888
rect 229706 162832 232116 162888
rect 229645 162830 232116 162832
rect 229645 162827 229711 162830
rect 353293 162210 353359 162213
rect 351900 162208 353359 162210
rect 351900 162152 353298 162208
rect 353354 162152 353359 162208
rect 351900 162150 353359 162152
rect 353293 162147 353359 162150
rect 229461 159082 229527 159085
rect 229461 159080 232116 159082
rect 229461 159024 229466 159080
rect 229522 159024 232116 159080
rect 229461 159022 232116 159024
rect 229461 159019 229527 159022
rect 353937 158674 354003 158677
rect 351900 158672 354003 158674
rect 351900 158616 353942 158672
rect 353998 158616 354003 158672
rect 351900 158614 354003 158616
rect 353937 158611 354003 158614
rect 230381 155274 230447 155277
rect 230381 155272 232116 155274
rect 230381 155216 230386 155272
rect 230442 155216 232116 155272
rect 230381 155214 232116 155216
rect 230381 155211 230447 155214
rect 353293 155138 353359 155141
rect 351900 155136 353359 155138
rect 351900 155080 353298 155136
rect 353354 155080 353359 155136
rect 351900 155078 353359 155080
rect 353293 155075 353359 155078
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 230381 151466 230447 151469
rect 353293 151466 353359 151469
rect 230381 151464 232116 151466
rect 230381 151408 230386 151464
rect 230442 151408 232116 151464
rect 230381 151406 232116 151408
rect 351900 151464 353359 151466
rect 351900 151408 353298 151464
rect 353354 151408 353359 151464
rect 351900 151406 353359 151408
rect 230381 151403 230447 151406
rect 353293 151403 353359 151406
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 354029 147930 354095 147933
rect 351900 147928 354095 147930
rect 351900 147872 354034 147928
rect 354090 147872 354095 147928
rect 351900 147870 354095 147872
rect 354029 147867 354095 147870
rect 229645 147658 229711 147661
rect 229645 147656 232116 147658
rect 229645 147600 229650 147656
rect 229706 147600 232116 147656
rect 229645 147598 232116 147600
rect 229645 147595 229711 147598
rect 353293 144394 353359 144397
rect 351900 144392 353359 144394
rect 351900 144336 353298 144392
rect 353354 144336 353359 144392
rect 351900 144334 353359 144336
rect 353293 144331 353359 144334
rect 230381 143850 230447 143853
rect 230381 143848 232116 143850
rect 230381 143792 230386 143848
rect 230442 143792 232116 143848
rect 230381 143790 232116 143792
rect 230381 143787 230447 143790
rect 353937 140858 354003 140861
rect 351900 140856 354003 140858
rect 351900 140800 353942 140856
rect 353998 140800 354003 140856
rect 351900 140798 354003 140800
rect 353937 140795 354003 140798
rect 230381 140042 230447 140045
rect 230381 140040 232116 140042
rect 230381 139984 230386 140040
rect 230442 139984 232116 140040
rect 230381 139982 232116 139984
rect 230381 139979 230447 139982
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 353293 137322 353359 137325
rect 351900 137320 353359 137322
rect 351900 137264 353298 137320
rect 353354 137264 353359 137320
rect 351900 137262 353359 137264
rect 353293 137259 353359 137262
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 229829 136234 229895 136237
rect 229829 136232 232116 136234
rect 229829 136176 229834 136232
rect 229890 136176 232116 136232
rect 229829 136174 232116 136176
rect 229829 136171 229895 136174
rect 354305 133786 354371 133789
rect 351900 133784 354371 133786
rect 351900 133728 354310 133784
rect 354366 133728 354371 133784
rect 351900 133726 354371 133728
rect 354305 133723 354371 133726
rect 229737 132426 229803 132429
rect 229737 132424 232116 132426
rect 229737 132368 229742 132424
rect 229798 132368 232116 132424
rect 229737 132366 232116 132368
rect 229737 132363 229803 132366
rect 353937 130250 354003 130253
rect 351900 130248 354003 130250
rect 351900 130192 353942 130248
rect 353998 130192 354003 130248
rect 351900 130190 354003 130192
rect 353937 130187 354003 130190
rect 230381 128618 230447 128621
rect 230381 128616 232116 128618
rect 230381 128560 230386 128616
rect 230442 128560 232116 128616
rect 230381 128558 232116 128560
rect 230381 128555 230447 128558
rect 354581 126578 354647 126581
rect 351900 126576 354647 126578
rect 351900 126520 354586 126576
rect 354642 126520 354647 126576
rect 351900 126518 354647 126520
rect 354581 126515 354647 126518
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 230105 124810 230171 124813
rect 230105 124808 232116 124810
rect 230105 124752 230110 124808
rect 230166 124752 232116 124808
rect 230105 124750 232116 124752
rect 230105 124747 230171 124750
rect -960 123572 480 123812
rect 354489 123042 354555 123045
rect 351900 123040 354555 123042
rect 351900 122984 354494 123040
rect 354550 122984 354555 123040
rect 351900 122982 354555 122984
rect 354489 122979 354555 122982
rect 230013 121002 230079 121005
rect 230013 121000 232116 121002
rect 230013 120944 230018 121000
rect 230074 120944 232116 121000
rect 230013 120942 232116 120944
rect 230013 120939 230079 120942
rect 354397 119506 354463 119509
rect 351900 119504 354463 119506
rect 351900 119448 354402 119504
rect 354458 119448 354463 119504
rect 351900 119446 354463 119448
rect 354397 119443 354463 119446
rect 230197 117194 230263 117197
rect 230197 117192 232116 117194
rect 230197 117136 230202 117192
rect 230258 117136 232116 117192
rect 230197 117134 232116 117136
rect 230197 117131 230263 117134
rect 354305 115970 354371 115973
rect 351900 115968 354371 115970
rect 351900 115912 354310 115968
rect 354366 115912 354371 115968
rect 351900 115910 354371 115912
rect 354305 115907 354371 115910
rect 229921 113386 229987 113389
rect 229921 113384 232116 113386
rect 229921 113328 229926 113384
rect 229982 113328 232116 113384
rect 229921 113326 232116 113328
rect 229921 113323 229987 113326
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 354213 112434 354279 112437
rect 351900 112432 354279 112434
rect 351900 112376 354218 112432
rect 354274 112376 354279 112432
rect 351900 112374 354279 112376
rect 354213 112371 354279 112374
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 229829 109578 229895 109581
rect 229829 109576 232116 109578
rect 229829 109520 229834 109576
rect 229890 109520 232116 109576
rect 229829 109518 232116 109520
rect 229829 109515 229895 109518
rect 354121 108898 354187 108901
rect 351900 108896 354187 108898
rect 351900 108840 354126 108896
rect 354182 108840 354187 108896
rect 351900 108838 354187 108840
rect 354121 108835 354187 108838
rect 230381 105770 230447 105773
rect 230381 105768 232116 105770
rect 230381 105712 230386 105768
rect 230442 105712 232116 105768
rect 230381 105710 232116 105712
rect 230381 105707 230447 105710
rect 354029 105362 354095 105365
rect 351900 105360 354095 105362
rect 351900 105304 354034 105360
rect 354090 105304 354095 105360
rect 351900 105302 354095 105304
rect 354029 105299 354095 105302
rect 229737 101962 229803 101965
rect 229737 101960 232116 101962
rect 229737 101904 229742 101960
rect 229798 101904 232116 101960
rect 229737 101902 232116 101904
rect 229737 101899 229803 101902
rect 353937 101826 354003 101829
rect 351900 101824 354003 101826
rect 351900 101768 353942 101824
rect 353998 101768 354003 101824
rect 351900 101766 354003 101768
rect 353937 101763 354003 101766
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 6453 3362 6519 3365
rect 233325 3362 233391 3365
rect 6453 3360 233391 3362
rect 6453 3304 6458 3360
rect 6514 3304 233330 3360
rect 233386 3304 233391 3360
rect 6453 3302 233391 3304
rect 6453 3299 6519 3302
rect 233325 3299 233391 3302
rect 351729 3362 351795 3365
rect 583385 3362 583451 3365
rect 351729 3360 583451 3362
rect 351729 3304 351734 3360
rect 351790 3304 583390 3360
rect 583446 3304 583451 3360
rect 351729 3302 583451 3304
rect 351729 3299 351795 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 262000 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 262000 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 262000 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 262000 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 262000 249914 286398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 262000 254414 290898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 262000 258914 295398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 262000 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 262000 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 262000 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 262000 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 262000 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 262000 285914 286398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 262000 290414 290898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 262000 294914 295398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 262000 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 262000 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 262000 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 262000 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 262000 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 262000 321914 286398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 262000 326414 290898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 262000 330914 295398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 262000 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 262000 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 262000 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 262000 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 262000 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 236208 255454 236528 255486
rect 236208 255218 236250 255454
rect 236486 255218 236528 255454
rect 236208 255134 236528 255218
rect 236208 254898 236250 255134
rect 236486 254898 236528 255134
rect 236208 254866 236528 254898
rect 266928 255454 267248 255486
rect 266928 255218 266970 255454
rect 267206 255218 267248 255454
rect 266928 255134 267248 255218
rect 266928 254898 266970 255134
rect 267206 254898 267248 255134
rect 266928 254866 267248 254898
rect 297648 255454 297968 255486
rect 297648 255218 297690 255454
rect 297926 255218 297968 255454
rect 297648 255134 297968 255218
rect 297648 254898 297690 255134
rect 297926 254898 297968 255134
rect 297648 254866 297968 254898
rect 328368 255454 328688 255486
rect 328368 255218 328410 255454
rect 328646 255218 328688 255454
rect 328368 255134 328688 255218
rect 328368 254898 328410 255134
rect 328646 254898 328688 255134
rect 328368 254866 328688 254898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 251568 223954 251888 223986
rect 251568 223718 251610 223954
rect 251846 223718 251888 223954
rect 251568 223634 251888 223718
rect 251568 223398 251610 223634
rect 251846 223398 251888 223634
rect 251568 223366 251888 223398
rect 282288 223954 282608 223986
rect 282288 223718 282330 223954
rect 282566 223718 282608 223954
rect 282288 223634 282608 223718
rect 282288 223398 282330 223634
rect 282566 223398 282608 223634
rect 282288 223366 282608 223398
rect 313008 223954 313328 223986
rect 313008 223718 313050 223954
rect 313286 223718 313328 223954
rect 313008 223634 313328 223718
rect 313008 223398 313050 223634
rect 313286 223398 313328 223634
rect 313008 223366 313328 223398
rect 343728 223954 344048 223986
rect 343728 223718 343770 223954
rect 344006 223718 344048 223954
rect 343728 223634 344048 223718
rect 343728 223398 343770 223634
rect 344006 223398 344048 223634
rect 343728 223366 344048 223398
rect 236208 219454 236528 219486
rect 236208 219218 236250 219454
rect 236486 219218 236528 219454
rect 236208 219134 236528 219218
rect 236208 218898 236250 219134
rect 236486 218898 236528 219134
rect 236208 218866 236528 218898
rect 266928 219454 267248 219486
rect 266928 219218 266970 219454
rect 267206 219218 267248 219454
rect 266928 219134 267248 219218
rect 266928 218898 266970 219134
rect 267206 218898 267248 219134
rect 266928 218866 267248 218898
rect 297648 219454 297968 219486
rect 297648 219218 297690 219454
rect 297926 219218 297968 219454
rect 297648 219134 297968 219218
rect 297648 218898 297690 219134
rect 297926 218898 297968 219134
rect 297648 218866 297968 218898
rect 328368 219454 328688 219486
rect 328368 219218 328410 219454
rect 328646 219218 328688 219454
rect 328368 219134 328688 219218
rect 328368 218898 328410 219134
rect 328646 218898 328688 219134
rect 328368 218866 328688 218898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 251568 187954 251888 187986
rect 251568 187718 251610 187954
rect 251846 187718 251888 187954
rect 251568 187634 251888 187718
rect 251568 187398 251610 187634
rect 251846 187398 251888 187634
rect 251568 187366 251888 187398
rect 282288 187954 282608 187986
rect 282288 187718 282330 187954
rect 282566 187718 282608 187954
rect 282288 187634 282608 187718
rect 282288 187398 282330 187634
rect 282566 187398 282608 187634
rect 282288 187366 282608 187398
rect 313008 187954 313328 187986
rect 313008 187718 313050 187954
rect 313286 187718 313328 187954
rect 313008 187634 313328 187718
rect 313008 187398 313050 187634
rect 313286 187398 313328 187634
rect 313008 187366 313328 187398
rect 343728 187954 344048 187986
rect 343728 187718 343770 187954
rect 344006 187718 344048 187954
rect 343728 187634 344048 187718
rect 343728 187398 343770 187634
rect 344006 187398 344048 187634
rect 343728 187366 344048 187398
rect 236208 183454 236528 183486
rect 236208 183218 236250 183454
rect 236486 183218 236528 183454
rect 236208 183134 236528 183218
rect 236208 182898 236250 183134
rect 236486 182898 236528 183134
rect 236208 182866 236528 182898
rect 266928 183454 267248 183486
rect 266928 183218 266970 183454
rect 267206 183218 267248 183454
rect 266928 183134 267248 183218
rect 266928 182898 266970 183134
rect 267206 182898 267248 183134
rect 266928 182866 267248 182898
rect 297648 183454 297968 183486
rect 297648 183218 297690 183454
rect 297926 183218 297968 183454
rect 297648 183134 297968 183218
rect 297648 182898 297690 183134
rect 297926 182898 297968 183134
rect 297648 182866 297968 182898
rect 328368 183454 328688 183486
rect 328368 183218 328410 183454
rect 328646 183218 328688 183454
rect 328368 183134 328688 183218
rect 328368 182898 328410 183134
rect 328646 182898 328688 183134
rect 328368 182866 328688 182898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 251568 151954 251888 151986
rect 251568 151718 251610 151954
rect 251846 151718 251888 151954
rect 251568 151634 251888 151718
rect 251568 151398 251610 151634
rect 251846 151398 251888 151634
rect 251568 151366 251888 151398
rect 282288 151954 282608 151986
rect 282288 151718 282330 151954
rect 282566 151718 282608 151954
rect 282288 151634 282608 151718
rect 282288 151398 282330 151634
rect 282566 151398 282608 151634
rect 282288 151366 282608 151398
rect 313008 151954 313328 151986
rect 313008 151718 313050 151954
rect 313286 151718 313328 151954
rect 313008 151634 313328 151718
rect 313008 151398 313050 151634
rect 313286 151398 313328 151634
rect 313008 151366 313328 151398
rect 343728 151954 344048 151986
rect 343728 151718 343770 151954
rect 344006 151718 344048 151954
rect 343728 151634 344048 151718
rect 343728 151398 343770 151634
rect 344006 151398 344048 151634
rect 343728 151366 344048 151398
rect 236208 147454 236528 147486
rect 236208 147218 236250 147454
rect 236486 147218 236528 147454
rect 236208 147134 236528 147218
rect 236208 146898 236250 147134
rect 236486 146898 236528 147134
rect 236208 146866 236528 146898
rect 266928 147454 267248 147486
rect 266928 147218 266970 147454
rect 267206 147218 267248 147454
rect 266928 147134 267248 147218
rect 266928 146898 266970 147134
rect 267206 146898 267248 147134
rect 266928 146866 267248 146898
rect 297648 147454 297968 147486
rect 297648 147218 297690 147454
rect 297926 147218 297968 147454
rect 297648 147134 297968 147218
rect 297648 146898 297690 147134
rect 297926 146898 297968 147134
rect 297648 146866 297968 146898
rect 328368 147454 328688 147486
rect 328368 147218 328410 147454
rect 328646 147218 328688 147454
rect 328368 147134 328688 147218
rect 328368 146898 328410 147134
rect 328646 146898 328688 147134
rect 328368 146866 328688 146898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 251568 115954 251888 115986
rect 251568 115718 251610 115954
rect 251846 115718 251888 115954
rect 251568 115634 251888 115718
rect 251568 115398 251610 115634
rect 251846 115398 251888 115634
rect 251568 115366 251888 115398
rect 282288 115954 282608 115986
rect 282288 115718 282330 115954
rect 282566 115718 282608 115954
rect 282288 115634 282608 115718
rect 282288 115398 282330 115634
rect 282566 115398 282608 115634
rect 282288 115366 282608 115398
rect 313008 115954 313328 115986
rect 313008 115718 313050 115954
rect 313286 115718 313328 115954
rect 313008 115634 313328 115718
rect 313008 115398 313050 115634
rect 313286 115398 313328 115634
rect 313008 115366 313328 115398
rect 343728 115954 344048 115986
rect 343728 115718 343770 115954
rect 344006 115718 344048 115954
rect 343728 115634 344048 115718
rect 343728 115398 343770 115634
rect 344006 115398 344048 115634
rect 343728 115366 344048 115398
rect 236208 111454 236528 111486
rect 236208 111218 236250 111454
rect 236486 111218 236528 111454
rect 236208 111134 236528 111218
rect 236208 110898 236250 111134
rect 236486 110898 236528 111134
rect 236208 110866 236528 110898
rect 266928 111454 267248 111486
rect 266928 111218 266970 111454
rect 267206 111218 267248 111454
rect 266928 111134 267248 111218
rect 266928 110898 266970 111134
rect 267206 110898 267248 111134
rect 266928 110866 267248 110898
rect 297648 111454 297968 111486
rect 297648 111218 297690 111454
rect 297926 111218 297968 111454
rect 297648 111134 297968 111218
rect 297648 110898 297690 111134
rect 297926 110898 297968 111134
rect 297648 110866 297968 110898
rect 328368 111454 328688 111486
rect 328368 111218 328410 111454
rect 328646 111218 328688 111454
rect 328368 111134 328688 111218
rect 328368 110898 328410 111134
rect 328646 110898 328688 111134
rect 328368 110866 328688 110898
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 88954 231914 98000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 98000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 97954 240914 98000
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 66454 245414 98000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 70954 249914 98000
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 75454 254414 98000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 79954 258914 98000
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 84454 263414 98000
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 88954 267914 98000
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 93454 272414 98000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 97954 276914 98000
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 66454 281414 98000
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 70954 285914 98000
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 75454 290414 98000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 79954 294914 98000
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 84454 299414 98000
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 88954 303914 98000
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 93454 308414 98000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 97954 312914 98000
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 98000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 70954 321914 98000
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 98000
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 79954 330914 98000
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 84454 335414 98000
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 88954 339914 98000
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 93454 344414 98000
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 97954 348914 98000
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 66454 353414 98000
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 236250 255218 236486 255454
rect 236250 254898 236486 255134
rect 266970 255218 267206 255454
rect 266970 254898 267206 255134
rect 297690 255218 297926 255454
rect 297690 254898 297926 255134
rect 328410 255218 328646 255454
rect 328410 254898 328646 255134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 251610 223718 251846 223954
rect 251610 223398 251846 223634
rect 282330 223718 282566 223954
rect 282330 223398 282566 223634
rect 313050 223718 313286 223954
rect 313050 223398 313286 223634
rect 343770 223718 344006 223954
rect 343770 223398 344006 223634
rect 236250 219218 236486 219454
rect 236250 218898 236486 219134
rect 266970 219218 267206 219454
rect 266970 218898 267206 219134
rect 297690 219218 297926 219454
rect 297690 218898 297926 219134
rect 328410 219218 328646 219454
rect 328410 218898 328646 219134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 251610 187718 251846 187954
rect 251610 187398 251846 187634
rect 282330 187718 282566 187954
rect 282330 187398 282566 187634
rect 313050 187718 313286 187954
rect 313050 187398 313286 187634
rect 343770 187718 344006 187954
rect 343770 187398 344006 187634
rect 236250 183218 236486 183454
rect 236250 182898 236486 183134
rect 266970 183218 267206 183454
rect 266970 182898 267206 183134
rect 297690 183218 297926 183454
rect 297690 182898 297926 183134
rect 328410 183218 328646 183454
rect 328410 182898 328646 183134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 251610 151718 251846 151954
rect 251610 151398 251846 151634
rect 282330 151718 282566 151954
rect 282330 151398 282566 151634
rect 313050 151718 313286 151954
rect 313050 151398 313286 151634
rect 343770 151718 344006 151954
rect 343770 151398 344006 151634
rect 236250 147218 236486 147454
rect 236250 146898 236486 147134
rect 266970 147218 267206 147454
rect 266970 146898 267206 147134
rect 297690 147218 297926 147454
rect 297690 146898 297926 147134
rect 328410 147218 328646 147454
rect 328410 146898 328646 147134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 251610 115718 251846 115954
rect 251610 115398 251846 115634
rect 282330 115718 282566 115954
rect 282330 115398 282566 115634
rect 313050 115718 313286 115954
rect 313050 115398 313286 115634
rect 343770 115718 344006 115954
rect 343770 115398 344006 115634
rect 236250 111218 236486 111454
rect 236250 110898 236486 111134
rect 266970 111218 267206 111454
rect 266970 110898 267206 111134
rect 297690 111218 297926 111454
rect 297690 110898 297926 111134
rect 328410 111218 328646 111454
rect 328410 110898 328646 111134
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 236250 255454
rect 236486 255218 266970 255454
rect 267206 255218 297690 255454
rect 297926 255218 328410 255454
rect 328646 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 236250 255134
rect 236486 254898 266970 255134
rect 267206 254898 297690 255134
rect 297926 254898 328410 255134
rect 328646 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 251610 223954
rect 251846 223718 282330 223954
rect 282566 223718 313050 223954
rect 313286 223718 343770 223954
rect 344006 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 251610 223634
rect 251846 223398 282330 223634
rect 282566 223398 313050 223634
rect 313286 223398 343770 223634
rect 344006 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 236250 219454
rect 236486 219218 266970 219454
rect 267206 219218 297690 219454
rect 297926 219218 328410 219454
rect 328646 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 236250 219134
rect 236486 218898 266970 219134
rect 267206 218898 297690 219134
rect 297926 218898 328410 219134
rect 328646 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 251610 187954
rect 251846 187718 282330 187954
rect 282566 187718 313050 187954
rect 313286 187718 343770 187954
rect 344006 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 251610 187634
rect 251846 187398 282330 187634
rect 282566 187398 313050 187634
rect 313286 187398 343770 187634
rect 344006 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 236250 183454
rect 236486 183218 266970 183454
rect 267206 183218 297690 183454
rect 297926 183218 328410 183454
rect 328646 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 236250 183134
rect 236486 182898 266970 183134
rect 267206 182898 297690 183134
rect 297926 182898 328410 183134
rect 328646 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 251610 151954
rect 251846 151718 282330 151954
rect 282566 151718 313050 151954
rect 313286 151718 343770 151954
rect 344006 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 251610 151634
rect 251846 151398 282330 151634
rect 282566 151398 313050 151634
rect 313286 151398 343770 151634
rect 344006 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 236250 147454
rect 236486 147218 266970 147454
rect 267206 147218 297690 147454
rect 297926 147218 328410 147454
rect 328646 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 236250 147134
rect 236486 146898 266970 147134
rect 267206 146898 297690 147134
rect 297926 146898 328410 147134
rect 328646 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 251610 115954
rect 251846 115718 282330 115954
rect 282566 115718 313050 115954
rect 313286 115718 343770 115954
rect 344006 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 251610 115634
rect 251846 115398 282330 115634
rect 282566 115398 313050 115634
rect 313286 115398 343770 115634
rect 344006 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 236250 111454
rect 236486 111218 266970 111454
rect 267206 111218 297690 111454
rect 297926 111218 328410 111454
rect 328646 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 236250 111134
rect 236486 110898 266970 111134
rect 267206 110898 297690 111134
rect 297926 110898 328410 111134
rect 328646 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 232000 0 1 100000
box 0 0 120000 160000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 98000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 262000 254414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 98000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 262000 290414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 98000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 262000 326414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 98000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 262000 263414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 98000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 262000 299414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 98000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 262000 335414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 98000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 262000 236414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 98000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 262000 272414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 98000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 262000 308414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 98000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 262000 344414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 98000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 262000 245414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 98000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 262000 281414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 98000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 262000 317414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 98000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 262000 353414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 98000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 262000 240914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 98000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 262000 276914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 98000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 262000 312914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 98000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 262000 348914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 98000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 262000 249914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 98000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 262000 285914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 98000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 262000 321914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 98000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 262000 258914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 98000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 262000 294914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 98000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 262000 330914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 98000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 262000 231914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 98000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 262000 267914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 98000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 262000 303914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 98000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 262000 339914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
