// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire \dff_last_analogFIGARO.D ;
 wire \dff_last_analogFIGARO.Q ;
 wire \dff_last_analogFIGARO.clk ;
 wire \dff_last_analogRO.D ;
 wire \dff_last_analogRO.Q ;
 wire \dff_last_sampledFIGARO.D ;
 wire \dff_last_sampledFIGARO.Q ;
 wire \dff_last_sampledRO.D ;
 wire \dff_last_sampledRO.Q ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[1] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[2] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[3] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[4] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[5] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[0] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[10] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[11] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[12] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[13] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[14] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[15] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[1] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[2] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[3] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[4] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[5] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[6] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[7] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[8] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[9] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[10] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[11] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[12] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[13] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[14] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[15] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[16] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[17] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[18] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[19] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[1] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[20] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[2] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[3] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[4] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[5] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[6] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[7] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[8] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[9] ;
 wire \entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ;
 wire \entropy_FIGARO.genblk1[1].dff_gen.Q ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[1] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[2] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[3] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[4] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[5] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[0] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[10] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[11] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[12] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[13] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[14] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[15] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[1] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[2] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[3] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[4] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[5] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[6] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[7] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[8] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[9] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[10] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[11] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[12] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[13] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[14] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[15] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[16] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[17] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[18] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[19] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[1] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[20] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[2] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[3] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[4] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[5] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[6] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[7] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[8] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[9] ;
 wire \entropy_FIGARO.genblk1[2].FIGARO_gen.o_figaro ;
 wire \entropy_FIGARO.genblk1[2].dff_gen.Q ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[1] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[2] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[3] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[4] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[5] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[0] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[10] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[11] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[12] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[13] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[14] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[15] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[1] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[2] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[3] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[4] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[5] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[6] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[7] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[8] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[9] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[10] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[11] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[12] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[13] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[14] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[15] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[16] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[17] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[18] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[19] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[1] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[20] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[2] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[3] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[4] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[5] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[6] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[7] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[8] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[9] ;
 wire \entropy_FIGARO.genblk1[3].FIGARO_gen.o_figaro ;
 wire \entropy_FIGARO.genblk1[3].dff_gen.Q ;
 wire \entropy_FIGARO.xor_stage.Xor_out[1] ;
 wire \entropy_FIGARO.xor_stage_analog.Xor_out[1] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[10].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[10].dff_gen.Q ;
 wire \entropy_RO.genblk1[11].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[11].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[11].dff_gen.Q ;
 wire \entropy_RO.genblk1[12].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[12].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[12].dff_gen.Q ;
 wire \entropy_RO.genblk1[13].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[13].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[13].dff_gen.Q ;
 wire \entropy_RO.genblk1[14].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[14].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[14].dff_gen.Q ;
 wire \entropy_RO.genblk1[15].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[15].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[15].dff_gen.Q ;
 wire \entropy_RO.genblk1[16].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[16].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[16].dff_gen.Q ;
 wire \entropy_RO.genblk1[17].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[17].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[17].dff_gen.Q ;
 wire \entropy_RO.genblk1[18].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[18].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[18].dff_gen.Q ;
 wire \entropy_RO.genblk1[19].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[19].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[19].dff_gen.Q ;
 wire \entropy_RO.genblk1[1].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[1].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[1].dff_gen.Q ;
 wire \entropy_RO.genblk1[20].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[20].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[20].dff_gen.Q ;
 wire \entropy_RO.genblk1[21].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[21].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[21].dff_gen.Q ;
 wire \entropy_RO.genblk1[22].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[22].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[22].dff_gen.Q ;
 wire \entropy_RO.genblk1[23].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[23].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[23].dff_gen.Q ;
 wire \entropy_RO.genblk1[24].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[24].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[24].dff_gen.Q ;
 wire \entropy_RO.genblk1[25].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[25].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[25].dff_gen.Q ;
 wire \entropy_RO.genblk1[26].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[26].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[26].dff_gen.Q ;
 wire \entropy_RO.genblk1[27].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[27].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[27].dff_gen.Q ;
 wire \entropy_RO.genblk1[28].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[28].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[28].dff_gen.Q ;
 wire \entropy_RO.genblk1[29].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[29].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[29].dff_gen.Q ;
 wire \entropy_RO.genblk1[2].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[2].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[2].dff_gen.Q ;
 wire \entropy_RO.genblk1[30].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[30].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[30].dff_gen.Q ;
 wire \entropy_RO.genblk1[31].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[31].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[31].dff_gen.Q ;
 wire \entropy_RO.genblk1[32].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[32].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[32].dff_gen.Q ;
 wire \entropy_RO.genblk1[33].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[33].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[33].dff_gen.Q ;
 wire \entropy_RO.genblk1[34].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[34].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[34].dff_gen.Q ;
 wire \entropy_RO.genblk1[35].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[35].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[35].dff_gen.Q ;
 wire \entropy_RO.genblk1[36].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[36].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[36].dff_gen.Q ;
 wire \entropy_RO.genblk1[37].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[37].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[37].dff_gen.Q ;
 wire \entropy_RO.genblk1[38].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[38].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[38].dff_gen.Q ;
 wire \entropy_RO.genblk1[39].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[39].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[39].dff_gen.Q ;
 wire \entropy_RO.genblk1[3].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[3].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[3].dff_gen.Q ;
 wire \entropy_RO.genblk1[40].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[40].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[40].dff_gen.Q ;
 wire \entropy_RO.genblk1[4].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[4].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[4].dff_gen.Q ;
 wire \entropy_RO.genblk1[5].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[5].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[5].dff_gen.Q ;
 wire \entropy_RO.genblk1[6].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[6].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[6].dff_gen.Q ;
 wire \entropy_RO.genblk1[7].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[7].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[7].dff_gen.Q ;
 wire \entropy_RO.genblk1[8].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[8].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[8].dff_gen.Q ;
 wire \entropy_RO.genblk1[9].RO_gen.del[0] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[10] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[11] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[12] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[13] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[14] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[1] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[2] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[3] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[4] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[5] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[6] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[7] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[8] ;
 wire \entropy_RO.genblk1[9].RO_gen.del[9] ;
 wire \entropy_RO.genblk1[9].dff_gen.Q ;
 wire \entropy_RO.xor_stage.Xor_out[10] ;
 wire \entropy_RO.xor_stage.Xor_out[11] ;
 wire \entropy_RO.xor_stage.Xor_out[12] ;
 wire \entropy_RO.xor_stage.Xor_out[13] ;
 wire \entropy_RO.xor_stage.Xor_out[14] ;
 wire \entropy_RO.xor_stage.Xor_out[15] ;
 wire \entropy_RO.xor_stage.Xor_out[16] ;
 wire \entropy_RO.xor_stage.Xor_out[17] ;
 wire \entropy_RO.xor_stage.Xor_out[18] ;
 wire \entropy_RO.xor_stage.Xor_out[19] ;
 wire \entropy_RO.xor_stage.Xor_out[1] ;
 wire \entropy_RO.xor_stage.Xor_out[20] ;
 wire \entropy_RO.xor_stage.Xor_out[21] ;
 wire \entropy_RO.xor_stage.Xor_out[22] ;
 wire \entropy_RO.xor_stage.Xor_out[23] ;
 wire \entropy_RO.xor_stage.Xor_out[24] ;
 wire \entropy_RO.xor_stage.Xor_out[25] ;
 wire \entropy_RO.xor_stage.Xor_out[26] ;
 wire \entropy_RO.xor_stage.Xor_out[27] ;
 wire \entropy_RO.xor_stage.Xor_out[28] ;
 wire \entropy_RO.xor_stage.Xor_out[29] ;
 wire \entropy_RO.xor_stage.Xor_out[2] ;
 wire \entropy_RO.xor_stage.Xor_out[30] ;
 wire \entropy_RO.xor_stage.Xor_out[31] ;
 wire \entropy_RO.xor_stage.Xor_out[32] ;
 wire \entropy_RO.xor_stage.Xor_out[33] ;
 wire \entropy_RO.xor_stage.Xor_out[34] ;
 wire \entropy_RO.xor_stage.Xor_out[35] ;
 wire \entropy_RO.xor_stage.Xor_out[36] ;
 wire \entropy_RO.xor_stage.Xor_out[37] ;
 wire \entropy_RO.xor_stage.Xor_out[38] ;
 wire \entropy_RO.xor_stage.Xor_out[3] ;
 wire \entropy_RO.xor_stage.Xor_out[4] ;
 wire \entropy_RO.xor_stage.Xor_out[5] ;
 wire \entropy_RO.xor_stage.Xor_out[6] ;
 wire \entropy_RO.xor_stage.Xor_out[7] ;
 wire \entropy_RO.xor_stage.Xor_out[8] ;
 wire \entropy_RO.xor_stage.Xor_out[9] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[10] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[11] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[12] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[13] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[14] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[15] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[16] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[17] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[18] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[19] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[1] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[20] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[21] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[22] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[23] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[24] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[25] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[26] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[27] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[28] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[29] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[2] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[30] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[31] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[32] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[33] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[34] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[35] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[36] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[37] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[38] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[3] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[4] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[5] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[6] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[7] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[8] ;
 wire \entropy_RO.xor_stage_analog.Xor_out[9] ;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire \clknet_0_dff_last_analogFIGARO.clk ;
 wire \clknet_1_0_0_dff_last_analogFIGARO.clk ;
 wire \clknet_1_0_1_dff_last_analogFIGARO.clk ;
 wire \clknet_1_1_0_dff_last_analogFIGARO.clk ;
 wire \clknet_1_1_1_dff_last_analogFIGARO.clk ;
 wire \clknet_2_0_0_dff_last_analogFIGARO.clk ;
 wire \clknet_2_0_1_dff_last_analogFIGARO.clk ;
 wire \clknet_2_1_0_dff_last_analogFIGARO.clk ;
 wire \clknet_2_1_1_dff_last_analogFIGARO.clk ;
 wire \clknet_2_2_0_dff_last_analogFIGARO.clk ;
 wire \clknet_2_2_1_dff_last_analogFIGARO.clk ;
 wire \clknet_2_3_0_dff_last_analogFIGARO.clk ;
 wire \clknet_2_3_1_dff_last_analogFIGARO.clk ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;

 sky130_fd_sc_hd__inv_2 _047_ (.A(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _048_ (.A(\dff_last_sampledRO.D ),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _049_ (.A(\dff_last_analogRO.D ),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _050_ (.A(\dff_last_sampledRO.Q ),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _051_ (.A(\dff_last_analogRO.Q ),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _052_ (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _053_ (.A(\dff_last_sampledFIGARO.D ),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _054_ (.A(\dff_last_analogFIGARO.D ),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _055_ (.A(\dff_last_sampledFIGARO.Q ),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _056_ (.A(\dff_last_analogFIGARO.Q ),
    .Y(_021_));
 sky130_fd_sc_hd__mux2_1 _057_ (.A0(la_data_in[64]),
    .A1(clknet_1_1__leaf_wb_clk_i),
    .S(la_oenb[64]),
    .X(\dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__and3b_2 _058_ (.A_N(wb_rst_i),
    .B(wbs_stb_i),
    .C(wbs_cyc_i),
    .X(_000_));
 sky130_fd_sc_hd__nand3b_2 _059_ (.A_N(wbs_we_i),
    .B(wbs_stb_i),
    .C(wbs_cyc_i),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_2 _060_ (.A(wbs_dat_o[6]),
    .B(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__or4_2 _061_ (.A(wbs_adr_i[5]),
    .B(wbs_adr_i[4]),
    .C(wbs_adr_i[7]),
    .D(wbs_adr_i[6]),
    .X(_024_));
 sky130_fd_sc_hd__or4b_2 _062_ (.A(wbs_adr_i[1]),
    .B(wbs_adr_i[0]),
    .C(wbs_adr_i[3]),
    .D_N(wbs_adr_i[2]),
    .X(_025_));
 sky130_fd_sc_hd__or4b_2 _063_ (.A(_022_),
    .B(_024_),
    .C(_025_),
    .D_N(net3),
    .X(_026_));
 sky130_fd_sc_hd__a21oi_2 _064_ (.A1(_023_),
    .A2(_026_),
    .B1(wb_rst_i),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_2 _065_ (.A(wbs_dat_o[1]),
    .B(_022_),
    .Y(_027_));
 sky130_fd_sc_hd__or4_2 _066_ (.A(_012_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_028_));
 sky130_fd_sc_hd__a21oi_2 _067_ (.A1(_027_),
    .A2(_028_),
    .B1(wb_rst_i),
    .Y(_002_));
 sky130_fd_sc_hd__nand2_2 _068_ (.A(wbs_dat_o[2]),
    .B(_022_),
    .Y(_029_));
 sky130_fd_sc_hd__or4_2 _069_ (.A(_013_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_030_));
 sky130_fd_sc_hd__a21oi_2 _070_ (.A1(_029_),
    .A2(_030_),
    .B1(wb_rst_i),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_2 _071_ (.A(wbs_dat_o[3]),
    .B(_022_),
    .Y(_031_));
 sky130_fd_sc_hd__or4_2 _072_ (.A(_014_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_032_));
 sky130_fd_sc_hd__a21oi_2 _073_ (.A1(_031_),
    .A2(_032_),
    .B1(wb_rst_i),
    .Y(_004_));
 sky130_fd_sc_hd__nand2_2 _074_ (.A(wbs_dat_o[4]),
    .B(_022_),
    .Y(_033_));
 sky130_fd_sc_hd__or4_2 _075_ (.A(_015_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_034_));
 sky130_fd_sc_hd__a21oi_2 _076_ (.A1(_033_),
    .A2(_034_),
    .B1(wb_rst_i),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_2 _077_ (.A(wbs_dat_o[5]),
    .B(_022_),
    .Y(_035_));
 sky130_fd_sc_hd__or4_2 _078_ (.A(_016_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_036_));
 sky130_fd_sc_hd__a21oi_2 _079_ (.A1(_035_),
    .A2(_036_),
    .B1(wb_rst_i),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_2 _080_ (.A(wbs_dat_o[7]),
    .B(_022_),
    .Y(_037_));
 sky130_fd_sc_hd__or4_2 _081_ (.A(_017_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_038_));
 sky130_fd_sc_hd__a21oi_2 _082_ (.A1(_037_),
    .A2(_038_),
    .B1(wb_rst_i),
    .Y(_007_));
 sky130_fd_sc_hd__nand2_2 _083_ (.A(wbs_dat_o[8]),
    .B(_022_),
    .Y(_039_));
 sky130_fd_sc_hd__or4_2 _084_ (.A(_018_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_040_));
 sky130_fd_sc_hd__a21oi_2 _085_ (.A1(_039_),
    .A2(_040_),
    .B1(wb_rst_i),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_2 _086_ (.A(wbs_dat_o[9]),
    .B(_022_),
    .Y(_041_));
 sky130_fd_sc_hd__or4_2 _087_ (.A(_019_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_042_));
 sky130_fd_sc_hd__a21oi_2 _088_ (.A1(_041_),
    .A2(_042_),
    .B1(wb_rst_i),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_2 _089_ (.A(wbs_dat_o[10]),
    .B(_022_),
    .Y(_043_));
 sky130_fd_sc_hd__or4_2 _090_ (.A(_020_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_044_));
 sky130_fd_sc_hd__a21oi_2 _091_ (.A1(_043_),
    .A2(_044_),
    .B1(wb_rst_i),
    .Y(_010_));
 sky130_fd_sc_hd__nand2_2 _092_ (.A(wbs_dat_o[11]),
    .B(_022_),
    .Y(_045_));
 sky130_fd_sc_hd__or4_2 _093_ (.A(_021_),
    .B(_022_),
    .C(_024_),
    .D(_025_),
    .X(_046_));
 sky130_fd_sc_hd__a21oi_2 _094_ (.A1(_045_),
    .A2(_046_),
    .B1(wb_rst_i),
    .Y(_011_));
 sky130_fd_sc_hd__dfxtp_2 _095_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_000_),
    .Q(wbs_ack_o));
 sky130_fd_sc_hd__dfxtp_2 _096_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_001_),
    .Q(wbs_dat_o[6]));
 sky130_fd_sc_hd__dfxtp_2 _097_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_002_),
    .Q(wbs_dat_o[1]));
 sky130_fd_sc_hd__dfxtp_2 _098_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_003_),
    .Q(wbs_dat_o[2]));
 sky130_fd_sc_hd__dfxtp_2 _099_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_004_),
    .Q(wbs_dat_o[3]));
 sky130_fd_sc_hd__dfxtp_2 _100_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_005_),
    .Q(wbs_dat_o[4]));
 sky130_fd_sc_hd__dfxtp_2 _101_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_006_),
    .Q(wbs_dat_o[5]));
 sky130_fd_sc_hd__dfxtp_2 _102_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_007_),
    .Q(wbs_dat_o[7]));
 sky130_fd_sc_hd__dfxtp_2 _103_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_008_),
    .Q(wbs_dat_o[8]));
 sky130_fd_sc_hd__dfxtp_2 _104_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_009_),
    .Q(wbs_dat_o[9]));
 sky130_fd_sc_hd__dfxtp_2 _105_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_010_),
    .Q(wbs_dat_o[10]));
 sky130_fd_sc_hd__dfxtp_2 _106_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_011_),
    .Q(wbs_dat_o[11]));
 sky130_fd_sc_hd__dfxtp_2 _107_ (.CLK(net12),
    .D(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[1].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _108_ (.CLK(net12),
    .D(\entropy_RO.genblk1[2].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[2].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _109_ (.CLK(net12),
    .D(\entropy_RO.genblk1[3].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[3].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _110_ (.CLK(net12),
    .D(\entropy_RO.genblk1[4].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[4].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _111_ (.CLK(net12),
    .D(\entropy_RO.genblk1[5].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[5].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _112_ (.CLK(net12),
    .D(\entropy_RO.genblk1[6].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[6].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _113_ (.CLK(net12),
    .D(\entropy_RO.genblk1[7].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[7].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _114_ (.CLK(\clknet_2_3_1_dff_last_analogFIGARO.clk ),
    .D(\entropy_RO.genblk1[8].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[8].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _115_ (.CLK(\clknet_2_3_1_dff_last_analogFIGARO.clk ),
    .D(\entropy_RO.genblk1[9].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[9].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _116_ (.CLK(\clknet_2_3_1_dff_last_analogFIGARO.clk ),
    .D(\entropy_RO.genblk1[10].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[10].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _117_ (.CLK(net15),
    .D(\entropy_RO.genblk1[11].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[11].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _118_ (.CLK(net15),
    .D(\entropy_RO.genblk1[12].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[12].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _119_ (.CLK(net15),
    .D(\entropy_RO.genblk1[13].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[13].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _120_ (.CLK(net15),
    .D(\entropy_RO.genblk1[14].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[14].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _121_ (.CLK(\clknet_2_1_1_dff_last_analogFIGARO.clk ),
    .D(\entropy_RO.genblk1[15].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[15].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _122_ (.CLK(net15),
    .D(\entropy_RO.genblk1[16].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[16].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _123_ (.CLK(net15),
    .D(\entropy_RO.genblk1[17].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[17].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _124_ (.CLK(net15),
    .D(\entropy_RO.genblk1[18].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[18].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _125_ (.CLK(net15),
    .D(\entropy_RO.genblk1[19].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[19].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _126_ (.CLK(net15),
    .D(\entropy_RO.genblk1[20].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[20].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _127_ (.CLK(net10),
    .D(\entropy_RO.genblk1[21].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[21].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _128_ (.CLK(net10),
    .D(\entropy_RO.genblk1[22].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[22].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _129_ (.CLK(net10),
    .D(\entropy_RO.genblk1[23].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[23].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _130_ (.CLK(net10),
    .D(\entropy_RO.genblk1[24].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[24].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _131_ (.CLK(net9),
    .D(\entropy_RO.genblk1[25].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[25].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _132_ (.CLK(net9),
    .D(\entropy_RO.genblk1[26].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[26].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _133_ (.CLK(net10),
    .D(\entropy_RO.genblk1[27].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[27].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _134_ (.CLK(net9),
    .D(\entropy_RO.genblk1[28].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[28].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _135_ (.CLK(net9),
    .D(\entropy_RO.genblk1[29].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[29].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _136_ (.CLK(net9),
    .D(\entropy_RO.genblk1[30].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[30].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _137_ (.CLK(net5),
    .D(\entropy_RO.genblk1[31].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[31].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _138_ (.CLK(net5),
    .D(\entropy_RO.genblk1[32].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[32].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _139_ (.CLK(net5),
    .D(\entropy_RO.genblk1[33].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[33].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _140_ (.CLK(net5),
    .D(\entropy_RO.genblk1[34].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[34].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _141_ (.CLK(net5),
    .D(\entropy_RO.genblk1[35].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[35].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _142_ (.CLK(net7),
    .D(\entropy_RO.genblk1[36].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[36].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _143_ (.CLK(net7),
    .D(\entropy_RO.genblk1[37].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[37].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _144_ (.CLK(net7),
    .D(\entropy_RO.genblk1[38].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[38].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _145_ (.CLK(net7),
    .D(\entropy_RO.genblk1[39].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[39].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _146_ (.CLK(net7),
    .D(\entropy_RO.genblk1[40].RO_gen.del[0] ),
    .Q(\entropy_RO.genblk1[40].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _147_ (.CLK(net4),
    .D(\dff_last_sampledRO.D ),
    .Q(\dff_last_sampledRO.Q ));
 sky130_fd_sc_hd__dfxtp_2 _148_ (.CLK(net3),
    .D(\dff_last_analogRO.D ),
    .Q(\dff_last_analogRO.Q ));
 sky130_fd_sc_hd__dfxtp_2 _149_ (.CLK(net9),
    .D(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ),
    .Q(\entropy_FIGARO.genblk1[1].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _150_ (.CLK(net9),
    .D(\entropy_FIGARO.genblk1[2].FIGARO_gen.o_figaro ),
    .Q(\entropy_FIGARO.genblk1[2].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _151_ (.CLK(net5),
    .D(\entropy_FIGARO.genblk1[3].FIGARO_gen.o_figaro ),
    .Q(\entropy_FIGARO.genblk1[3].dff_gen.Q ));
 sky130_fd_sc_hd__dfxtp_2 _152_ (.CLK(net11),
    .D(\dff_last_sampledFIGARO.D ),
    .Q(\dff_last_sampledFIGARO.Q ));
 sky130_fd_sc_hd__dfxtp_2 _153_ (.CLK(net11),
    .D(\dff_last_analogFIGARO.D ),
    .Q(\dff_last_analogFIGARO.Q ));
 sky130_fd_sc_hd__conb_1 _154_ (.HI(io_oeb[0]));
 sky130_fd_sc_hd__conb_1 _155_ (.HI(io_oeb[1]));
 sky130_fd_sc_hd__conb_1 _156_ (.HI(io_oeb[2]));
 sky130_fd_sc_hd__conb_1 _157_ (.HI(io_oeb[3]));
 sky130_fd_sc_hd__conb_1 _158_ (.HI(io_oeb[4]));
 sky130_fd_sc_hd__conb_1 _159_ (.HI(io_oeb[5]));
 sky130_fd_sc_hd__conb_1 _160_ (.HI(io_oeb[6]));
 sky130_fd_sc_hd__conb_1 _161_ (.HI(io_oeb[7]));
 sky130_fd_sc_hd__conb_1 _162_ (.HI(io_oeb[8]));
 sky130_fd_sc_hd__conb_1 _163_ (.HI(io_oeb[9]));
 sky130_fd_sc_hd__conb_1 _164_ (.HI(io_oeb[10]));
 sky130_fd_sc_hd__conb_1 _165_ (.HI(io_oeb[11]));
 sky130_fd_sc_hd__conb_1 _166_ (.HI(io_oeb[12]));
 sky130_fd_sc_hd__conb_1 _167_ (.HI(io_oeb[13]));
 sky130_fd_sc_hd__conb_1 _168_ (.HI(io_oeb[14]));
 sky130_fd_sc_hd__conb_1 _169_ (.HI(io_oeb[15]));
 sky130_fd_sc_hd__conb_1 _170_ (.HI(io_oeb[16]));
 sky130_fd_sc_hd__conb_1 _171_ (.HI(io_oeb[17]));
 sky130_fd_sc_hd__conb_1 _172_ (.HI(io_oeb[18]));
 sky130_fd_sc_hd__conb_1 _173_ (.HI(io_oeb[19]));
 sky130_fd_sc_hd__conb_1 _174_ (.HI(io_oeb[20]));
 sky130_fd_sc_hd__conb_1 _175_ (.HI(io_oeb[21]));
 sky130_fd_sc_hd__conb_1 _176_ (.HI(io_oeb[22]));
 sky130_fd_sc_hd__conb_1 _177_ (.HI(io_oeb[23]));
 sky130_fd_sc_hd__conb_1 _178_ (.HI(io_oeb[24]));
 sky130_fd_sc_hd__conb_1 _179_ (.HI(io_oeb[25]));
 sky130_fd_sc_hd__conb_1 _180_ (.HI(io_oeb[26]));
 sky130_fd_sc_hd__conb_1 _181_ (.HI(io_oeb[27]));
 sky130_fd_sc_hd__conb_1 _182_ (.HI(io_oeb[28]));
 sky130_fd_sc_hd__conb_1 _183_ (.HI(io_oeb[29]));
 sky130_fd_sc_hd__conb_1 _184_ (.HI(io_oeb[30]));
 sky130_fd_sc_hd__conb_1 _185_ (.HI(io_oeb[31]));
 sky130_fd_sc_hd__conb_1 _186_ (.HI(io_oeb[32]));
 sky130_fd_sc_hd__conb_1 _187_ (.HI(io_oeb[33]));
 sky130_fd_sc_hd__conb_1 _188_ (.HI(io_oeb[34]));
 sky130_fd_sc_hd__conb_1 _189_ (.HI(io_oeb[35]));
 sky130_fd_sc_hd__conb_1 _190_ (.HI(io_oeb[36]));
 sky130_fd_sc_hd__conb_1 _191_ (.LO(io_oeb[37]));
 sky130_fd_sc_hd__conb_1 _192_ (.LO(io_out[12]));
 sky130_fd_sc_hd__conb_1 _193_ (.LO(io_out[13]));
 sky130_fd_sc_hd__conb_1 _194_ (.LO(io_out[14]));
 sky130_fd_sc_hd__conb_1 _195_ (.LO(io_out[15]));
 sky130_fd_sc_hd__conb_1 _196_ (.LO(io_out[16]));
 sky130_fd_sc_hd__conb_1 _197_ (.LO(io_out[17]));
 sky130_fd_sc_hd__conb_1 _198_ (.LO(io_out[18]));
 sky130_fd_sc_hd__conb_1 _199_ (.LO(io_out[19]));
 sky130_fd_sc_hd__conb_1 _200_ (.LO(io_out[32]));
 sky130_fd_sc_hd__conb_1 _201_ (.LO(io_out[33]));
 sky130_fd_sc_hd__conb_1 _202_ (.LO(io_out[34]));
 sky130_fd_sc_hd__conb_1 _203_ (.LO(io_out[35]));
 sky130_fd_sc_hd__conb_1 _204_ (.LO(io_out[36]));
 sky130_fd_sc_hd__conb_1 _205_ (.LO(io_out[37]));
 sky130_fd_sc_hd__conb_1 _206_ (.LO(irq[0]));
 sky130_fd_sc_hd__conb_1 _207_ (.LO(irq[1]));
 sky130_fd_sc_hd__conb_1 _208_ (.LO(irq[2]));
 sky130_fd_sc_hd__conb_1 _209_ (.LO(la_data_out[12]));
 sky130_fd_sc_hd__conb_1 _210_ (.LO(la_data_out[13]));
 sky130_fd_sc_hd__conb_1 _211_ (.LO(la_data_out[14]));
 sky130_fd_sc_hd__conb_1 _212_ (.LO(la_data_out[15]));
 sky130_fd_sc_hd__conb_1 _213_ (.LO(la_data_out[16]));
 sky130_fd_sc_hd__conb_1 _214_ (.LO(la_data_out[17]));
 sky130_fd_sc_hd__conb_1 _215_ (.LO(la_data_out[18]));
 sky130_fd_sc_hd__conb_1 _216_ (.LO(la_data_out[19]));
 sky130_fd_sc_hd__conb_1 _217_ (.LO(la_data_out[20]));
 sky130_fd_sc_hd__conb_1 _218_ (.LO(la_data_out[21]));
 sky130_fd_sc_hd__conb_1 _219_ (.LO(la_data_out[22]));
 sky130_fd_sc_hd__conb_1 _220_ (.LO(la_data_out[23]));
 sky130_fd_sc_hd__conb_1 _221_ (.LO(la_data_out[24]));
 sky130_fd_sc_hd__conb_1 _222_ (.LO(la_data_out[25]));
 sky130_fd_sc_hd__conb_1 _223_ (.LO(la_data_out[26]));
 sky130_fd_sc_hd__conb_1 _224_ (.LO(la_data_out[27]));
 sky130_fd_sc_hd__conb_1 _225_ (.LO(la_data_out[28]));
 sky130_fd_sc_hd__conb_1 _226_ (.LO(la_data_out[29]));
 sky130_fd_sc_hd__conb_1 _227_ (.LO(la_data_out[30]));
 sky130_fd_sc_hd__conb_1 _228_ (.LO(la_data_out[31]));
 sky130_fd_sc_hd__conb_1 _229_ (.LO(la_data_out[44]));
 sky130_fd_sc_hd__conb_1 _230_ (.LO(la_data_out[45]));
 sky130_fd_sc_hd__conb_1 _231_ (.LO(la_data_out[46]));
 sky130_fd_sc_hd__conb_1 _232_ (.LO(la_data_out[47]));
 sky130_fd_sc_hd__conb_1 _233_ (.LO(la_data_out[48]));
 sky130_fd_sc_hd__conb_1 _234_ (.LO(la_data_out[49]));
 sky130_fd_sc_hd__conb_1 _235_ (.LO(la_data_out[50]));
 sky130_fd_sc_hd__conb_1 _236_ (.LO(la_data_out[51]));
 sky130_fd_sc_hd__conb_1 _237_ (.LO(la_data_out[52]));
 sky130_fd_sc_hd__conb_1 _238_ (.LO(la_data_out[53]));
 sky130_fd_sc_hd__conb_1 _239_ (.LO(la_data_out[54]));
 sky130_fd_sc_hd__conb_1 _240_ (.LO(la_data_out[55]));
 sky130_fd_sc_hd__conb_1 _241_ (.LO(la_data_out[56]));
 sky130_fd_sc_hd__conb_1 _242_ (.LO(la_data_out[57]));
 sky130_fd_sc_hd__conb_1 _243_ (.LO(la_data_out[58]));
 sky130_fd_sc_hd__conb_1 _244_ (.LO(la_data_out[59]));
 sky130_fd_sc_hd__conb_1 _245_ (.LO(la_data_out[60]));
 sky130_fd_sc_hd__conb_1 _246_ (.LO(la_data_out[61]));
 sky130_fd_sc_hd__conb_1 _247_ (.LO(la_data_out[62]));
 sky130_fd_sc_hd__conb_1 _248_ (.LO(la_data_out[63]));
 sky130_fd_sc_hd__conb_1 _249_ (.LO(la_data_out[64]));
 sky130_fd_sc_hd__conb_1 _250_ (.LO(la_data_out[65]));
 sky130_fd_sc_hd__conb_1 _251_ (.LO(la_data_out[66]));
 sky130_fd_sc_hd__conb_1 _252_ (.LO(la_data_out[67]));
 sky130_fd_sc_hd__conb_1 _253_ (.LO(la_data_out[68]));
 sky130_fd_sc_hd__conb_1 _254_ (.LO(la_data_out[69]));
 sky130_fd_sc_hd__conb_1 _255_ (.LO(la_data_out[70]));
 sky130_fd_sc_hd__conb_1 _256_ (.LO(la_data_out[71]));
 sky130_fd_sc_hd__conb_1 _257_ (.LO(la_data_out[72]));
 sky130_fd_sc_hd__conb_1 _258_ (.LO(la_data_out[73]));
 sky130_fd_sc_hd__conb_1 _259_ (.LO(la_data_out[74]));
 sky130_fd_sc_hd__conb_1 _260_ (.LO(la_data_out[75]));
 sky130_fd_sc_hd__conb_1 _261_ (.LO(la_data_out[76]));
 sky130_fd_sc_hd__conb_1 _262_ (.LO(la_data_out[77]));
 sky130_fd_sc_hd__conb_1 _263_ (.LO(la_data_out[78]));
 sky130_fd_sc_hd__conb_1 _264_ (.LO(la_data_out[79]));
 sky130_fd_sc_hd__conb_1 _265_ (.LO(la_data_out[80]));
 sky130_fd_sc_hd__conb_1 _266_ (.LO(la_data_out[81]));
 sky130_fd_sc_hd__conb_1 _267_ (.LO(la_data_out[82]));
 sky130_fd_sc_hd__conb_1 _268_ (.LO(la_data_out[83]));
 sky130_fd_sc_hd__conb_1 _269_ (.LO(la_data_out[84]));
 sky130_fd_sc_hd__conb_1 _270_ (.LO(la_data_out[85]));
 sky130_fd_sc_hd__conb_1 _271_ (.LO(la_data_out[86]));
 sky130_fd_sc_hd__conb_1 _272_ (.LO(la_data_out[87]));
 sky130_fd_sc_hd__conb_1 _273_ (.LO(la_data_out[88]));
 sky130_fd_sc_hd__conb_1 _274_ (.LO(la_data_out[89]));
 sky130_fd_sc_hd__conb_1 _275_ (.LO(la_data_out[90]));
 sky130_fd_sc_hd__conb_1 _276_ (.LO(la_data_out[91]));
 sky130_fd_sc_hd__conb_1 _277_ (.LO(la_data_out[92]));
 sky130_fd_sc_hd__conb_1 _278_ (.LO(la_data_out[93]));
 sky130_fd_sc_hd__conb_1 _279_ (.LO(la_data_out[94]));
 sky130_fd_sc_hd__conb_1 _280_ (.LO(la_data_out[95]));
 sky130_fd_sc_hd__conb_1 _281_ (.LO(la_data_out[96]));
 sky130_fd_sc_hd__conb_1 _282_ (.LO(la_data_out[97]));
 sky130_fd_sc_hd__conb_1 _283_ (.LO(la_data_out[98]));
 sky130_fd_sc_hd__conb_1 _284_ (.LO(la_data_out[99]));
 sky130_fd_sc_hd__conb_1 _285_ (.LO(la_data_out[100]));
 sky130_fd_sc_hd__conb_1 _286_ (.LO(la_data_out[101]));
 sky130_fd_sc_hd__conb_1 _287_ (.LO(la_data_out[102]));
 sky130_fd_sc_hd__conb_1 _288_ (.LO(la_data_out[103]));
 sky130_fd_sc_hd__conb_1 _289_ (.LO(la_data_out[104]));
 sky130_fd_sc_hd__conb_1 _290_ (.LO(la_data_out[105]));
 sky130_fd_sc_hd__conb_1 _291_ (.LO(la_data_out[106]));
 sky130_fd_sc_hd__conb_1 _292_ (.LO(la_data_out[107]));
 sky130_fd_sc_hd__conb_1 _293_ (.LO(la_data_out[108]));
 sky130_fd_sc_hd__conb_1 _294_ (.LO(la_data_out[109]));
 sky130_fd_sc_hd__conb_1 _295_ (.LO(la_data_out[110]));
 sky130_fd_sc_hd__conb_1 _296_ (.LO(la_data_out[111]));
 sky130_fd_sc_hd__conb_1 _297_ (.LO(la_data_out[112]));
 sky130_fd_sc_hd__conb_1 _298_ (.LO(la_data_out[113]));
 sky130_fd_sc_hd__conb_1 _299_ (.LO(la_data_out[114]));
 sky130_fd_sc_hd__conb_1 _300_ (.LO(la_data_out[115]));
 sky130_fd_sc_hd__conb_1 _301_ (.LO(la_data_out[116]));
 sky130_fd_sc_hd__conb_1 _302_ (.LO(la_data_out[117]));
 sky130_fd_sc_hd__conb_1 _303_ (.LO(la_data_out[118]));
 sky130_fd_sc_hd__conb_1 _304_ (.LO(la_data_out[119]));
 sky130_fd_sc_hd__conb_1 _305_ (.LO(la_data_out[120]));
 sky130_fd_sc_hd__conb_1 _306_ (.LO(la_data_out[121]));
 sky130_fd_sc_hd__conb_1 _307_ (.LO(la_data_out[122]));
 sky130_fd_sc_hd__conb_1 _308_ (.LO(la_data_out[123]));
 sky130_fd_sc_hd__conb_1 _309_ (.LO(la_data_out[124]));
 sky130_fd_sc_hd__conb_1 _310_ (.LO(la_data_out[125]));
 sky130_fd_sc_hd__conb_1 _311_ (.LO(la_data_out[126]));
 sky130_fd_sc_hd__conb_1 _312_ (.LO(la_data_out[127]));
 sky130_fd_sc_hd__conb_1 _313_ (.LO(wbs_dat_o[12]));
 sky130_fd_sc_hd__conb_1 _314_ (.LO(wbs_dat_o[13]));
 sky130_fd_sc_hd__conb_1 _315_ (.LO(wbs_dat_o[14]));
 sky130_fd_sc_hd__conb_1 _316_ (.LO(wbs_dat_o[15]));
 sky130_fd_sc_hd__conb_1 _317_ (.LO(wbs_dat_o[16]));
 sky130_fd_sc_hd__conb_1 _318_ (.LO(wbs_dat_o[17]));
 sky130_fd_sc_hd__conb_1 _319_ (.LO(wbs_dat_o[18]));
 sky130_fd_sc_hd__conb_1 _320_ (.LO(wbs_dat_o[19]));
 sky130_fd_sc_hd__conb_1 _321_ (.LO(wbs_dat_o[20]));
 sky130_fd_sc_hd__conb_1 _322_ (.LO(wbs_dat_o[21]));
 sky130_fd_sc_hd__conb_1 _323_ (.LO(wbs_dat_o[22]));
 sky130_fd_sc_hd__conb_1 _324_ (.LO(wbs_dat_o[23]));
 sky130_fd_sc_hd__conb_1 _325_ (.LO(wbs_dat_o[24]));
 sky130_fd_sc_hd__conb_1 _326_ (.LO(wbs_dat_o[25]));
 sky130_fd_sc_hd__conb_1 _327_ (.LO(wbs_dat_o[26]));
 sky130_fd_sc_hd__conb_1 _328_ (.LO(wbs_dat_o[27]));
 sky130_fd_sc_hd__conb_1 _329_ (.LO(wbs_dat_o[28]));
 sky130_fd_sc_hd__conb_1 _330_ (.LO(wbs_dat_o[29]));
 sky130_fd_sc_hd__conb_1 _331_ (.LO(wbs_dat_o[30]));
 sky130_fd_sc_hd__conb_1 _332_ (.LO(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_4 _333_ (.A(net6),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 _334_ (.A(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 _335_ (.A(\dff_last_sampledRO.D ),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 _336_ (.A(\dff_last_analogRO.D ),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 _337_ (.A(\dff_last_sampledRO.Q ),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 _338_ (.A(\dff_last_analogRO.Q ),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 _339_ (.A(net8),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 _340_ (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_4 _341_ (.A(\dff_last_sampledFIGARO.D ),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_4 _342_ (.A(\dff_last_analogFIGARO.D ),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_4 _343_ (.A(\dff_last_sampledFIGARO.Q ),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_4 _344_ (.A(\dff_last_analogFIGARO.Q ),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_4 _345_ (.A(net13),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 _346_ (.A(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 _347_ (.A(\dff_last_sampledRO.D ),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_4 _348_ (.A(\dff_last_analogRO.D ),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_4 _349_ (.A(\dff_last_sampledRO.Q ),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_4 _350_ (.A(\dff_last_analogRO.Q ),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_4 _351_ (.A(net11),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_4 _352_ (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_4 _353_ (.A(\dff_last_sampledFIGARO.D ),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_4 _354_ (.A(\dff_last_analogFIGARO.D ),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_4 _355_ (.A(\dff_last_sampledFIGARO.Q ),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_4 _356_ (.A(\dff_last_analogFIGARO.Q ),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_4 _357_ (.A(net4),
    .X(la_data_out[0]));
 sky130_fd_sc_hd__buf_4 _358_ (.A(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .X(la_data_out[1]));
 sky130_fd_sc_hd__buf_4 _359_ (.A(\dff_last_sampledRO.D ),
    .X(la_data_out[2]));
 sky130_fd_sc_hd__buf_4 _360_ (.A(\dff_last_analogRO.D ),
    .X(la_data_out[3]));
 sky130_fd_sc_hd__buf_4 _361_ (.A(\dff_last_sampledRO.Q ),
    .X(la_data_out[4]));
 sky130_fd_sc_hd__buf_4 _362_ (.A(\dff_last_analogRO.Q ),
    .X(la_data_out[5]));
 sky130_fd_sc_hd__buf_4 _363_ (.A(net4),
    .X(la_data_out[6]));
 sky130_fd_sc_hd__buf_4 _364_ (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ),
    .X(la_data_out[7]));
 sky130_fd_sc_hd__buf_4 _365_ (.A(\dff_last_sampledFIGARO.D ),
    .X(la_data_out[8]));
 sky130_fd_sc_hd__buf_4 _366_ (.A(\dff_last_analogFIGARO.D ),
    .X(la_data_out[9]));
 sky130_fd_sc_hd__buf_4 _367_ (.A(\dff_last_sampledFIGARO.Q ),
    .X(la_data_out[10]));
 sky130_fd_sc_hd__buf_4 _368_ (.A(\dff_last_analogFIGARO.Q ),
    .X(la_data_out[11]));
 sky130_fd_sc_hd__buf_4 _369_ (.A(net4),
    .X(la_data_out[32]));
 sky130_fd_sc_hd__buf_4 _370_ (.A(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .X(la_data_out[33]));
 sky130_fd_sc_hd__buf_4 _371_ (.A(\dff_last_sampledRO.D ),
    .X(la_data_out[34]));
 sky130_fd_sc_hd__buf_4 _372_ (.A(\dff_last_analogRO.D ),
    .X(la_data_out[35]));
 sky130_fd_sc_hd__buf_4 _373_ (.A(\dff_last_sampledRO.Q ),
    .X(la_data_out[36]));
 sky130_fd_sc_hd__buf_4 _374_ (.A(\dff_last_analogRO.Q ),
    .X(la_data_out[37]));
 sky130_fd_sc_hd__buf_4 _375_ (.A(net4),
    .X(la_data_out[38]));
 sky130_fd_sc_hd__buf_4 _376_ (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ),
    .X(la_data_out[39]));
 sky130_fd_sc_hd__buf_4 _377_ (.A(\dff_last_sampledFIGARO.D ),
    .X(la_data_out[40]));
 sky130_fd_sc_hd__buf_4 _378_ (.A(\dff_last_analogFIGARO.D ),
    .X(la_data_out[41]));
 sky130_fd_sc_hd__buf_4 _379_ (.A(\dff_last_sampledFIGARO.Q ),
    .X(la_data_out[42]));
 sky130_fd_sc_hd__buf_4 _380_ (.A(\dff_last_analogFIGARO.Q ),
    .X(la_data_out[43]));
 sky130_fd_sc_hd__buf_4 _381_ (.A(wbs_dat_o[6]),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[0].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[0] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[10].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[10] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[11].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[11] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[12].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[12] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[13].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[13] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[14].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[14] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[15] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[1].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[1] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[2].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[2] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[3].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[3] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[4].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[4] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[5].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[5] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[6].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[6] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[7].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[7] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[8].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[8] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.genblk1[9].inverters  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[9] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[10] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.xor_firo_1  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[15] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[14] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.xor_firo_2  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[5] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[7] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[4] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.xor_firo_3  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[4] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[6] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[3] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.xor_firo_4  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[3] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[5] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.xor_firo_5  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[2] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[4] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[1] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.firo.xor_firo_6  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.fXor[1] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[2] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter1  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[1] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter10  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[15] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter11  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[16] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[15] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter12  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[17] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[16] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter13  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[18] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[17] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter14  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[19] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[18] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter15  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[20] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter2  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[2] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter3  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[4] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter4  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[5] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter5  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[7] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter6  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[9] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter7  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[11] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter8  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[13] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.inverter9  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[14] ),
    .Y(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[13] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.xor_garo_1  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[3] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.xor_garo_2  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[6] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.xor_garo_3  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[8] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[7] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.xor_garo_4  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[10] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[9] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.xor_garo_5  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[12] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[11] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.garo.xor_garo_6  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[20] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[19] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[1].FIGARO_gen.xor_poly3  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[1].FIGARO_gen.firo.f[15] ),
    .X(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[0].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[0] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[10].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[10] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[11].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[11] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[12].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[12] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[13].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[13] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[14].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[14] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[15] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[1].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[1] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[2].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[2] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[3].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[3] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[4].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[4] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[5].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[5] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[6].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[6] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[7].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[7] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[8].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[8] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.genblk1[9].inverters  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[9] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[10] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.xor_firo_1  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[15] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[14] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.xor_firo_2  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[5] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[7] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[4] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.xor_firo_3  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[4] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[6] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[3] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.xor_firo_4  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[3] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[5] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.xor_firo_5  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[2] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[4] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[1] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.firo.xor_firo_6  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.fXor[1] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[2] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter1  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[1] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter10  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[15] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter11  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[16] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[15] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter12  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[17] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[16] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter13  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[18] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[17] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter14  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[19] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[18] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter15  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[20] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter2  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[2] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter3  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[4] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter4  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[5] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter5  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[7] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter6  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[9] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter7  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[11] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter8  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[13] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.inverter9  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[14] ),
    .Y(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[13] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.xor_garo_1  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[3] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.xor_garo_2  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[6] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.xor_garo_3  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[8] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[7] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.xor_garo_4  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[10] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[9] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.xor_garo_5  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[12] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[11] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.garo.xor_garo_6  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[20] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[19] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[2].FIGARO_gen.xor_poly3  (.A(\entropy_FIGARO.genblk1[2].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.firo.f[15] ),
    .X(\entropy_FIGARO.genblk1[2].FIGARO_gen.o_figaro ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[0].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[0] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[10].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[10] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[11].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[11] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[12].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[12] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[13].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[13] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[14].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[14] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[15] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[1].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[1] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[2].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[2] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[3].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[3] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[4].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[4] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[5].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[5] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[6].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[6] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[7].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[7] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[8].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[8] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.genblk1[9].inverters  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[9] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[10] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.xor_firo_1  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[15] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[14] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.xor_firo_2  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[5] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[7] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[4] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.xor_firo_3  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[4] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[6] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[3] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.xor_firo_4  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[3] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[5] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.xor_firo_5  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[2] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[4] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[1] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.firo.xor_firo_6  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.fXor[1] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[2] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter1  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[1] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter10  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[15] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter11  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[16] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[15] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter12  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[17] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[16] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter13  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[18] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[17] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter14  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[19] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[18] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter15  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[20] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter2  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[2] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter3  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[4] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter4  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[5] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter5  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[7] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter6  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[9] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter7  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[11] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter8  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[13] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.inverter9  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[14] ),
    .Y(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[13] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.xor_garo_1  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[3] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.xor_garo_2  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[6] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.xor_garo_3  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[8] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[7] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.xor_garo_4  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[10] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[9] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.xor_garo_5  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[12] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[11] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.garo.xor_garo_6  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[20] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[19] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.genblk1[3].FIGARO_gen.xor_poly3  (.A(\entropy_FIGARO.genblk1[3].FIGARO_gen.garo.f[0] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.firo.f[15] ),
    .X(\entropy_FIGARO.genblk1[3].FIGARO_gen.o_figaro ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.xor_stage.genblk1[1].xors  (.A(\entropy_FIGARO.xor_stage.Xor_out[1] ),
    .B(\entropy_FIGARO.genblk1[3].dff_gen.Q ),
    .X(\dff_last_analogFIGARO.D ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.xor_stage.xor_initial  (.A(\entropy_FIGARO.genblk1[1].dff_gen.Q ),
    .B(\entropy_FIGARO.genblk1[2].dff_gen.Q ),
    .X(\entropy_FIGARO.xor_stage.Xor_out[1] ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.xor_stage_analog.genblk1[1].xors  (.A(\entropy_FIGARO.xor_stage_analog.Xor_out[1] ),
    .B(\entropy_FIGARO.genblk1[3].FIGARO_gen.o_figaro ),
    .X(\dff_last_sampledFIGARO.D ));
 sky130_fd_sc_hd__xor2_4 \entropy_FIGARO.xor_stage_analog.xor_initial  (.A(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ),
    .B(\entropy_FIGARO.genblk1[2].FIGARO_gen.o_figaro ),
    .X(\entropy_FIGARO.xor_stage_analog.Xor_out[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[10].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[10].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[10].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[11].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[11].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[11].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[12].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[12].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[12].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[13].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[13].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[13].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[14].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[14].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[14].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[15].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[15].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[15].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[16].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[16].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[16].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[17].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[17].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[17].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[18].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[18].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[18].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[19].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[19].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[19].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[1].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[1].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[1].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[20].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[20].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[20].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[21].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[21].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[21].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[22].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[22].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[22].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[23].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[23].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[23].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[24].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[24].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[24].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[25].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[25].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[25].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[26].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[26].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[26].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[27].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[27].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[27].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[28].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[28].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[28].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[29].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[29].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[29].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[2].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[2].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[2].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[30].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[30].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[30].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[31].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[31].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[31].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[32].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[32].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[32].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[33].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[33].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[33].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[34].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[34].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[34].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[35].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[35].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[35].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[36].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[36].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[36].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[37].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[37].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[37].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[38].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[38].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[38].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[39].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[39].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[39].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[3].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[3].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[3].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[40].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[40].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[40].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[4].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[4].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[4].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[5].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[5].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[5].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[6].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[6].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[6].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[7].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[7].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[7].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[8].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[8].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[8].RO_gen.del[10] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[0].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[0] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[1] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[10].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[10] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[11] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[11].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[11] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[12] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[12].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[12] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[13] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[13].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[13] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[14] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[14].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[14] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[0] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[1].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[1] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[2] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[2].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[2] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[3] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[3].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[3] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[4] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[4].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[4] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[5] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[5].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[5] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[6] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[6].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[6] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[7] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[7].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[7] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[8] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[8].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[8] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[9] ));
 sky130_fd_sc_hd__inv_2 \entropy_RO.genblk1[9].RO_gen.genblk1[9].inverters  (.A(\entropy_RO.genblk1[9].RO_gen.del[9] ),
    .Y(\entropy_RO.genblk1[9].RO_gen.del[10] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[10].xors  (.A(\entropy_RO.xor_stage.Xor_out[10] ),
    .B(\entropy_RO.genblk1[12].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[11] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[11].xors  (.A(\entropy_RO.xor_stage.Xor_out[11] ),
    .B(\entropy_RO.genblk1[13].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[12] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[12].xors  (.A(\entropy_RO.xor_stage.Xor_out[12] ),
    .B(\entropy_RO.genblk1[14].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[13] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[13].xors  (.A(\entropy_RO.xor_stage.Xor_out[13] ),
    .B(\entropy_RO.genblk1[15].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[14] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[14].xors  (.A(\entropy_RO.xor_stage.Xor_out[14] ),
    .B(\entropy_RO.genblk1[16].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[15] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[15].xors  (.A(\entropy_RO.xor_stage.Xor_out[15] ),
    .B(\entropy_RO.genblk1[17].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[16] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[16].xors  (.A(\entropy_RO.xor_stage.Xor_out[16] ),
    .B(\entropy_RO.genblk1[18].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[17] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[17].xors  (.A(\entropy_RO.xor_stage.Xor_out[17] ),
    .B(\entropy_RO.genblk1[19].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[18] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[18].xors  (.A(\entropy_RO.xor_stage.Xor_out[18] ),
    .B(\entropy_RO.genblk1[20].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[19] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[19].xors  (.A(\entropy_RO.xor_stage.Xor_out[19] ),
    .B(\entropy_RO.genblk1[21].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[20] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[1].xors  (.A(\entropy_RO.xor_stage.Xor_out[1] ),
    .B(\entropy_RO.genblk1[3].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[20].xors  (.A(\entropy_RO.xor_stage.Xor_out[20] ),
    .B(\entropy_RO.genblk1[22].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[21] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[21].xors  (.A(\entropy_RO.xor_stage.Xor_out[21] ),
    .B(\entropy_RO.genblk1[23].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[22] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[22].xors  (.A(\entropy_RO.xor_stage.Xor_out[22] ),
    .B(\entropy_RO.genblk1[24].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[23] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[23].xors  (.A(\entropy_RO.xor_stage.Xor_out[23] ),
    .B(\entropy_RO.genblk1[25].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[24] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[24].xors  (.A(\entropy_RO.xor_stage.Xor_out[24] ),
    .B(\entropy_RO.genblk1[26].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[25] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[25].xors  (.A(\entropy_RO.xor_stage.Xor_out[25] ),
    .B(\entropy_RO.genblk1[27].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[26] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[26].xors  (.A(\entropy_RO.xor_stage.Xor_out[26] ),
    .B(\entropy_RO.genblk1[28].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[27] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[27].xors  (.A(\entropy_RO.xor_stage.Xor_out[27] ),
    .B(\entropy_RO.genblk1[29].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[28] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[28].xors  (.A(\entropy_RO.xor_stage.Xor_out[28] ),
    .B(\entropy_RO.genblk1[30].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[29] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[29].xors  (.A(\entropy_RO.xor_stage.Xor_out[29] ),
    .B(\entropy_RO.genblk1[31].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[30] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[2].xors  (.A(\entropy_RO.xor_stage.Xor_out[2] ),
    .B(\entropy_RO.genblk1[4].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[3] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[30].xors  (.A(\entropy_RO.xor_stage.Xor_out[30] ),
    .B(\entropy_RO.genblk1[32].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[31] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[31].xors  (.A(\entropy_RO.xor_stage.Xor_out[31] ),
    .B(\entropy_RO.genblk1[33].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[32] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[32].xors  (.A(\entropy_RO.xor_stage.Xor_out[32] ),
    .B(\entropy_RO.genblk1[34].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[33] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[33].xors  (.A(\entropy_RO.xor_stage.Xor_out[33] ),
    .B(\entropy_RO.genblk1[35].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[34] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[34].xors  (.A(\entropy_RO.xor_stage.Xor_out[34] ),
    .B(\entropy_RO.genblk1[36].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[35] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[35].xors  (.A(\entropy_RO.xor_stage.Xor_out[35] ),
    .B(\entropy_RO.genblk1[37].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[36] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[36].xors  (.A(\entropy_RO.xor_stage.Xor_out[36] ),
    .B(\entropy_RO.genblk1[38].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[37] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[37].xors  (.A(\entropy_RO.xor_stage.Xor_out[37] ),
    .B(\entropy_RO.genblk1[39].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[38] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[38].xors  (.A(\entropy_RO.xor_stage.Xor_out[38] ),
    .B(\entropy_RO.genblk1[40].dff_gen.Q ),
    .X(\dff_last_sampledRO.D ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[3].xors  (.A(\entropy_RO.xor_stage.Xor_out[3] ),
    .B(\entropy_RO.genblk1[5].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[4] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[4].xors  (.A(\entropy_RO.xor_stage.Xor_out[4] ),
    .B(\entropy_RO.genblk1[6].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[5].xors  (.A(\entropy_RO.xor_stage.Xor_out[5] ),
    .B(\entropy_RO.genblk1[7].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[6] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[6].xors  (.A(\entropy_RO.xor_stage.Xor_out[6] ),
    .B(\entropy_RO.genblk1[8].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[7] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[7].xors  (.A(\entropy_RO.xor_stage.Xor_out[7] ),
    .B(\entropy_RO.genblk1[9].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[8] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[8].xors  (.A(\entropy_RO.xor_stage.Xor_out[8] ),
    .B(\entropy_RO.genblk1[10].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[9] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.genblk1[9].xors  (.A(\entropy_RO.xor_stage.Xor_out[9] ),
    .B(\entropy_RO.genblk1[11].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[10] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage.xor_initial  (.A(\entropy_RO.genblk1[1].dff_gen.Q ),
    .B(\entropy_RO.genblk1[2].dff_gen.Q ),
    .X(\entropy_RO.xor_stage.Xor_out[1] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[10].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[10] ),
    .B(\entropy_RO.genblk1[12].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[11] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[11].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[11] ),
    .B(\entropy_RO.genblk1[13].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[12] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[12].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[12] ),
    .B(\entropy_RO.genblk1[14].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[13] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[13].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[13] ),
    .B(\entropy_RO.genblk1[15].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[14] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[14].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[14] ),
    .B(\entropy_RO.genblk1[16].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[15] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[15].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[15] ),
    .B(\entropy_RO.genblk1[17].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[16] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[16].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[16] ),
    .B(\entropy_RO.genblk1[18].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[17] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[17].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[17] ),
    .B(\entropy_RO.genblk1[19].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[18] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[18].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[18] ),
    .B(\entropy_RO.genblk1[20].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[19] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[19].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[19] ),
    .B(\entropy_RO.genblk1[21].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[20] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[1].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[1] ),
    .B(\entropy_RO.genblk1[3].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[2] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[20].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[20] ),
    .B(\entropy_RO.genblk1[22].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[21] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[21].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[21] ),
    .B(\entropy_RO.genblk1[23].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[22] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[22].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[22] ),
    .B(\entropy_RO.genblk1[24].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[23] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[23].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[23] ),
    .B(\entropy_RO.genblk1[25].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[24] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[24].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[24] ),
    .B(\entropy_RO.genblk1[26].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[25] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[25].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[25] ),
    .B(\entropy_RO.genblk1[27].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[26] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[26].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[26] ),
    .B(\entropy_RO.genblk1[28].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[27] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[27].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[27] ),
    .B(\entropy_RO.genblk1[29].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[28] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[28].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[28] ),
    .B(\entropy_RO.genblk1[30].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[29] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[29].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[29] ),
    .B(\entropy_RO.genblk1[31].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[30] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[2].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[2] ),
    .B(\entropy_RO.genblk1[4].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[3] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[30].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[30] ),
    .B(\entropy_RO.genblk1[32].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[31] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[31].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[31] ),
    .B(\entropy_RO.genblk1[33].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[32] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[32].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[32] ),
    .B(\entropy_RO.genblk1[34].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[33] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[33].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[33] ),
    .B(\entropy_RO.genblk1[35].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[34] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[34].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[34] ),
    .B(\entropy_RO.genblk1[36].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[35] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[35].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[35] ),
    .B(\entropy_RO.genblk1[37].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[36] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[36].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[36] ),
    .B(\entropy_RO.genblk1[38].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[37] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[37].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[37] ),
    .B(\entropy_RO.genblk1[39].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[38] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[38].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[38] ),
    .B(\entropy_RO.genblk1[40].RO_gen.del[0] ),
    .X(\dff_last_analogRO.D ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[3].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[3] ),
    .B(\entropy_RO.genblk1[5].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[4] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[4].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[4] ),
    .B(\entropy_RO.genblk1[6].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[5] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[5].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[5] ),
    .B(\entropy_RO.genblk1[7].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[6] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[6].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[6] ),
    .B(\entropy_RO.genblk1[8].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[7] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[7].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[7] ),
    .B(\entropy_RO.genblk1[9].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[8] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[8].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[8] ),
    .B(\entropy_RO.genblk1[10].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[9] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.genblk1[9].xors  (.A(\entropy_RO.xor_stage_analog.Xor_out[9] ),
    .B(\entropy_RO.genblk1[11].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[10] ));
 sky130_fd_sc_hd__xor2_4 \entropy_RO.xor_stage_analog.xor_initial  (.A(\entropy_RO.genblk1[1].RO_gen.del[0] ),
    .B(\entropy_RO.genblk1[2].RO_gen.del[0] ),
    .X(\entropy_RO.xor_stage_analog.Xor_out[1] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dff_last_analogFIGARO.clk  (.A(net1),
    .X(\clknet_0_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_0_0_dff_last_analogFIGARO.clk  (.A(\clknet_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_1_0_0_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_0_1_dff_last_analogFIGARO.clk  (.A(\clknet_1_0_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_1_0_1_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_1_0_dff_last_analogFIGARO.clk  (.A(\clknet_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_1_1_0_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_1_1_dff_last_analogFIGARO.clk  (.A(\clknet_1_1_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_1_1_1_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_0_0_dff_last_analogFIGARO.clk  (.A(\clknet_1_0_1_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_0_0_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_0_1_dff_last_analogFIGARO.clk  (.A(\clknet_2_0_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_0_1_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_1_0_dff_last_analogFIGARO.clk  (.A(\clknet_1_0_1_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_1_0_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_1_1_dff_last_analogFIGARO.clk  (.A(\clknet_2_1_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_1_1_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_2_0_dff_last_analogFIGARO.clk  (.A(\clknet_1_1_1_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_2_0_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_2_1_dff_last_analogFIGARO.clk  (.A(\clknet_2_2_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_2_1_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_3_0_dff_last_analogFIGARO.clk  (.A(\clknet_1_1_1_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_3_0_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_3_1_dff_last_analogFIGARO.clk  (.A(\clknet_2_3_0_dff_last_analogFIGARO.clk ),
    .X(\clknet_2_3_1_dff_last_analogFIGARO.clk ));
 sky130_fd_sc_hd__buf_4 wire1 (.A(net2),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 wire2 (.A(\dff_last_analogFIGARO.clk ),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 wire3 (.A(net4),
    .X(net3));
 sky130_fd_sc_hd__buf_2 wire4 (.A(\clknet_2_0_1_dff_last_analogFIGARO.clk ),
    .X(net4));
 sky130_fd_sc_hd__buf_2 max_length5 (.A(net7),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 wire6 (.A(net7),
    .X(net6));
 sky130_fd_sc_hd__buf_2 wire7 (.A(\clknet_2_0_1_dff_last_analogFIGARO.clk ),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 wire8 (.A(\clknet_2_1_1_dff_last_analogFIGARO.clk ),
    .X(net8));
 sky130_fd_sc_hd__buf_2 max_length9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_length10 (.A(\clknet_2_1_1_dff_last_analogFIGARO.clk ),
    .X(net10));
 sky130_fd_sc_hd__buf_2 wire11 (.A(\clknet_2_2_1_dff_last_analogFIGARO.clk ),
    .X(net11));
 sky130_fd_sc_hd__buf_2 wire12 (.A(\clknet_2_2_1_dff_last_analogFIGARO.clk ),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 wire13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 wire14 (.A(\clknet_2_3_1_dff_last_analogFIGARO.clk ),
    .X(net14));
 sky130_fd_sc_hd__buf_2 max_length15 (.A(\clknet_2_3_1_dff_last_analogFIGARO.clk ),
    .X(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\dff_last_analogFIGARO.D ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\dff_last_analogRO.D ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\dff_last_analogRO.D ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\dff_last_sampledFIGARO.D ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\dff_last_sampledFIGARO.D ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\dff_last_sampledRO.D ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\entropy_FIGARO.genblk1[1].FIGARO_gen.o_figaro ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(la_oenb[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net11));
 sky130_fd_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_355 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_360 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_158 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_317 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_334 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_369 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_526 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_598 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_610 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_730 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_773 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_777 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_831 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_848 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_875 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_890 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_954 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1000 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1111 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1122 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1146 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_239 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1127 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1136 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1148 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1172 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_339 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_427 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_431 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_443 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_512 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_565 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_880 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_892 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_916 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_955 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1101 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1118 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1124 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1136 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_241 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_274 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_158 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_227 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_620 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_632 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1276 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_187 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_199 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_238 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_244 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_256 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_268 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_355 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_367 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_273 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_217 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_240 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_272 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_273 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_179 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_248 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_272 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_160 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_194 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_255 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_834 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_776 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_819 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_831 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_843 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_775 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_819 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_831 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_843 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_988 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1000 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1012 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1024 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_750 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_832 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_774 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_866 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_722 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_793 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_847 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_856 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_868 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_892 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_716 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_728 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_845 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_866 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_704 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_847 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_859 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_871 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_833 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_842 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_625 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_637 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_760 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_772 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_636 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_636 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_648 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_660 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_719 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_833 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_838 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_862 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_688 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_719 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_731 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_850 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_862 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_894 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_705 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_723 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_216 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_694 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_703 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_754 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_778 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_676 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_679 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_696 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_666 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_777 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_782 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_806 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_625 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_637 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_750 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_681 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_721 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_679 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_688 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_700 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_762 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_694 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_750 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_668 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_747 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_782 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_829 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_722 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_76 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_692 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_719 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_731 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_788 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_591 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_542 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_603 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_651 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_694 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_471 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_679 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_688 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_700 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_724 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_653 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_677 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_694 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_569 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_524 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_580 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_511 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_523 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_535 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_691 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_700 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_724 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_488 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_500 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_524 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_719 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_731 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_720 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_715 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_777 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_786 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_610 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_690 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_483 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_495 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_582 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_790 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_496 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_612 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_483 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_495 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_547 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_582 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_709 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_778 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_469 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_651 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_663 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_675 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_726 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_750 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_469 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_474 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_498 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_520 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_532 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_556 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_649 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_677 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_700 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_724 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_576 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_660 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_511 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_523 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_535 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_579 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_679 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_691 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_703 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_507 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_659 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_663 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_675 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_788 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_787 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_808 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_647 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_693 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_776 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_539 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_543 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_555 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_607 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_651 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_663 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_675 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_726 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_750 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_776 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_788 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_554 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_648 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_720 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_660 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_721 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_744 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_579 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_604 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_664 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_675 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_567 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_579 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_591 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_649 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_680 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_692 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_704 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_716 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_632 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_722 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_627 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_636 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_648 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_660 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_735 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_747 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_759 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_540 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_549 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_651 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_663 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_675 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_724 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_102_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_539 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_548 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_639 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_648 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_660 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_735 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_747 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_759 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_103_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_593 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_660 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_104_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_105_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_486 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_498 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_566 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_106_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_458 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_500 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_792 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_804 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_816 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_828 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_107_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_502 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_526 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_788 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_108_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_455 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_467 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_498 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_626 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_638 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_109_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_435 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_444 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_468 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_110_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_511 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_523 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_535 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_698 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_722 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_111_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_434 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_443 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_526 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_112_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_511 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_523 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_535 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_621 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_625 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_637 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_113_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_114_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_115_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_610 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_619 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_661 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_116_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_624 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_666 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_117_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_622 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_625 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_612 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_636 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_121_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_625 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_627 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_649 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_667 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_718 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_630 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_639 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_735 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_747 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_759 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_125_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_638 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_719 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_728 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_647 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_720 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_778 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_127_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_607 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_611 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_786 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_812 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_836 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_129_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_665 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_779 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_788 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_130_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_647 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_131_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_694 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_765 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_132_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_632 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_644 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_668 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_737 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_756 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_780 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_133_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_619 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_640 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_134_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_135_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_609 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_618 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_136_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_666 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_137_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_726 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_782 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_806 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_138_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_698 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_722 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_139_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_651 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_646 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_690 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_749 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_772 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_141_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_520 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_721 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_786 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_142_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_469 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_520 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_567 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_579 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_689 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_698 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_812 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_836 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_143_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_560 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_523 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_567 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_576 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_588 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_612 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_633 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_679 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_683 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_695 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_812 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_836 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_145_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_582 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_786 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_810 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_146_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_526 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_567 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_579 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_591 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_147_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_524 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_552 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_754 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_778 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_719 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_776 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_812 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_836 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_151_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_497 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_520 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_800 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_152_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_17 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_153_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_484 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_496 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_508 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_520 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_582 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_777 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_786 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_154_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_155_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_488 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_497 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_597 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_721 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_156_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_523 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_554 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_610 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_681 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_157_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_427 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_439 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_490 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_499 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_558 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_582 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_705 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_728 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_765 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_770 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_782 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_806 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_440 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_481 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_513 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_679 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_776 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_159_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_443 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_452 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_464 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_677 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_722 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_772 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_160_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_444 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_525 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_637 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_791 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_803 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_815 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_161_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_442 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_772 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_162_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_355 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_367 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_163_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_584 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_164_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_608 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_687 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_165_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_556 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_653 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_166_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_567 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_576 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_588 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_612 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_722 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_167_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_271 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_555 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_564 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_576 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_719 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_728 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_168_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_735 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_747 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_759 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_169_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_734 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_170_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_469 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_586 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_668 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_735 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_744 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_756 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_780 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_171_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_621 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_730 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_172_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_639 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_695 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_704 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_735 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_747 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_759 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_173_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_716 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_728 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_174_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_175_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_707 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_716 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_728 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_752 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_176_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_40 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_700 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_177_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_626 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_638 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_179_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_180_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_301 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_181_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_182_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_183_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_184_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_185_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_186_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_187_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_189_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_190_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_21 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_191_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_192_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_9 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_17 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_193_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_194_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_195_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_196_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_197_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_198_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_199_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_200_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_201_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_202_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_203_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_204_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_205_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_206_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_207_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_209_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_210_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_211_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_212_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_213_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_214_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_215_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_216_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_217_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_218_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_219_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_220_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_221_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_222_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_223_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_224_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_225_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_226_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_583 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_227_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_228_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_229_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_230_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_231_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_232_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_233_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_234_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_235_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_236_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_17 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_237_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_238_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_239_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_240_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_241_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_242_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_243_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_244_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_245_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_246_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_247_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_248_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_249_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_250_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_251_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_252_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_253_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_254_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_255_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_256_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_257_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_258_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_259_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_260_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_261_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_262_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_263_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_264_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_265_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_266_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_267_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_268_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_269_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_270_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_271_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_272_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_273_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_274_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_275_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_276_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_277_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_278_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_279_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_280_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_281_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_194 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_450 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_474 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_498 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_530 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_595 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_607 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_733 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_750 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_877 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_882 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_894 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_931 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_943 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_955 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_1034 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_1069 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1086 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1168 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1180 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_1213 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1218 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1230 ();
 sky130_fd_sc_hd__decap_12 FILLER_282_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_1275 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_615 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_685 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_727 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_741 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_783 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_797 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_839 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_853 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_895 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_909 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_951 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_965 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1007 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1021 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1063 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1077 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1119 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1133 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1175 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1189 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1231 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1245 ();
 sky130_fd_sc_hd__decap_12 FILLER_283_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_1269 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_657 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_699 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_713 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_769 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_811 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_825 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_867 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_881 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_923 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_937 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_979 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_993 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1035 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1049 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1091 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1105 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1147 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1161 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1203 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1217 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1259 ();
 sky130_fd_sc_hd__decap_12 FILLER_284_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_1273 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_669 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_697 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_701 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_725 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_729 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_753 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_757 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_781 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_785 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_809 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_813 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_837 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_841 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_865 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_869 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_893 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_897 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_921 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_925 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_949 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_953 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_977 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_981 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1005 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1009 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1033 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1037 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1061 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1065 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1089 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1093 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1117 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1121 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1145 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1149 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1173 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1177 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1201 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1205 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1229 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1233 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1257 ();
 sky130_fd_sc_hd__decap_12 FILLER_285_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_1273 ();
endmodule

