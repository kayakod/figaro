magic
tech sky130B
magscale 1 2
timestamp 1669988164
<< obsli1 >>
rect 1104 2159 118864 157777
<< obsm1 >>
rect 1104 2128 118864 157808
<< metal2 >>
rect 2502 159200 2558 160000
rect 6918 159200 6974 160000
rect 11334 159200 11390 160000
rect 15750 159200 15806 160000
rect 20166 159200 20222 160000
rect 24582 159200 24638 160000
rect 28998 159200 29054 160000
rect 33414 159200 33470 160000
rect 37830 159200 37886 160000
rect 42246 159200 42302 160000
rect 46662 159200 46718 160000
rect 51078 159200 51134 160000
rect 55494 159200 55550 160000
rect 59910 159200 59966 160000
rect 64326 159200 64382 160000
rect 68742 159200 68798 160000
rect 73158 159200 73214 160000
rect 77574 159200 77630 160000
rect 81990 159200 82046 160000
rect 86406 159200 86462 160000
rect 90822 159200 90878 160000
rect 95238 159200 95294 160000
rect 99654 159200 99710 160000
rect 104070 159200 104126 160000
rect 108486 159200 108542 160000
rect 112902 159200 112958 160000
rect 117318 159200 117374 160000
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79230 0 79286 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90638 0 90694 800
rect 90822 0 90878 800
rect 91006 0 91062 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92478 0 92534 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94686 0 94742 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96158 0 96214 800
rect 96342 0 96398 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98182 0 98238 800
rect 98366 0 98422 800
rect 98550 0 98606 800
rect 98734 0 98790 800
rect 98918 0 98974 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
rect 100022 0 100078 800
rect 100206 0 100262 800
rect 100390 0 100446 800
rect 100574 0 100630 800
rect 100758 0 100814 800
rect 100942 0 100998 800
rect 101126 0 101182 800
rect 101310 0 101366 800
rect 101494 0 101550 800
rect 101678 0 101734 800
rect 101862 0 101918 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102414 0 102470 800
rect 102598 0 102654 800
rect 102782 0 102838 800
rect 102966 0 103022 800
rect 103150 0 103206 800
rect 103334 0 103390 800
rect 103518 0 103574 800
rect 103702 0 103758 800
rect 103886 0 103942 800
rect 104070 0 104126 800
rect 104254 0 104310 800
rect 104438 0 104494 800
rect 104622 0 104678 800
rect 104806 0 104862 800
rect 104990 0 105046 800
rect 105174 0 105230 800
<< obsm2 >>
rect 2136 159144 2446 159338
rect 2614 159144 6862 159338
rect 7030 159144 11278 159338
rect 11446 159144 15694 159338
rect 15862 159144 20110 159338
rect 20278 159144 24526 159338
rect 24694 159144 28942 159338
rect 29110 159144 33358 159338
rect 33526 159144 37774 159338
rect 37942 159144 42190 159338
rect 42358 159144 46606 159338
rect 46774 159144 51022 159338
rect 51190 159144 55438 159338
rect 55606 159144 59854 159338
rect 60022 159144 64270 159338
rect 64438 159144 68686 159338
rect 68854 159144 73102 159338
rect 73270 159144 77518 159338
rect 77686 159144 81934 159338
rect 82102 159144 86350 159338
rect 86518 159144 90766 159338
rect 90934 159144 95182 159338
rect 95350 159144 99598 159338
rect 99766 159144 104014 159338
rect 104182 159144 108430 159338
rect 108598 159144 112846 159338
rect 113014 159144 117262 159338
rect 117430 159144 117742 159338
rect 2136 856 117742 159144
rect 2136 800 14590 856
rect 14758 800 14774 856
rect 14942 800 14958 856
rect 15126 800 15142 856
rect 15310 800 15326 856
rect 15494 800 15510 856
rect 15678 800 15694 856
rect 15862 800 15878 856
rect 16046 800 16062 856
rect 16230 800 16246 856
rect 16414 800 16430 856
rect 16598 800 16614 856
rect 16782 800 16798 856
rect 16966 800 16982 856
rect 17150 800 17166 856
rect 17334 800 17350 856
rect 17518 800 17534 856
rect 17702 800 17718 856
rect 17886 800 17902 856
rect 18070 800 18086 856
rect 18254 800 18270 856
rect 18438 800 18454 856
rect 18622 800 18638 856
rect 18806 800 18822 856
rect 18990 800 19006 856
rect 19174 800 19190 856
rect 19358 800 19374 856
rect 19542 800 19558 856
rect 19726 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20110 856
rect 20278 800 20294 856
rect 20462 800 20478 856
rect 20646 800 20662 856
rect 20830 800 20846 856
rect 21014 800 21030 856
rect 21198 800 21214 856
rect 21382 800 21398 856
rect 21566 800 21582 856
rect 21750 800 21766 856
rect 21934 800 21950 856
rect 22118 800 22134 856
rect 22302 800 22318 856
rect 22486 800 22502 856
rect 22670 800 22686 856
rect 22854 800 22870 856
rect 23038 800 23054 856
rect 23222 800 23238 856
rect 23406 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23790 856
rect 23958 800 23974 856
rect 24142 800 24158 856
rect 24326 800 24342 856
rect 24510 800 24526 856
rect 24694 800 24710 856
rect 24878 800 24894 856
rect 25062 800 25078 856
rect 25246 800 25262 856
rect 25430 800 25446 856
rect 25614 800 25630 856
rect 25798 800 25814 856
rect 25982 800 25998 856
rect 26166 800 26182 856
rect 26350 800 26366 856
rect 26534 800 26550 856
rect 26718 800 26734 856
rect 26902 800 26918 856
rect 27086 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27654 856
rect 27822 800 27838 856
rect 28006 800 28022 856
rect 28190 800 28206 856
rect 28374 800 28390 856
rect 28558 800 28574 856
rect 28742 800 28758 856
rect 28926 800 28942 856
rect 29110 800 29126 856
rect 29294 800 29310 856
rect 29478 800 29494 856
rect 29662 800 29678 856
rect 29846 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30230 856
rect 30398 800 30414 856
rect 30582 800 30598 856
rect 30766 800 30782 856
rect 30950 800 30966 856
rect 31134 800 31150 856
rect 31318 800 31334 856
rect 31502 800 31518 856
rect 31686 800 31702 856
rect 31870 800 31886 856
rect 32054 800 32070 856
rect 32238 800 32254 856
rect 32422 800 32438 856
rect 32606 800 32622 856
rect 32790 800 32806 856
rect 32974 800 32990 856
rect 33158 800 33174 856
rect 33342 800 33358 856
rect 33526 800 33542 856
rect 33710 800 33726 856
rect 33894 800 33910 856
rect 34078 800 34094 856
rect 34262 800 34278 856
rect 34446 800 34462 856
rect 34630 800 34646 856
rect 34814 800 34830 856
rect 34998 800 35014 856
rect 35182 800 35198 856
rect 35366 800 35382 856
rect 35550 800 35566 856
rect 35734 800 35750 856
rect 35918 800 35934 856
rect 36102 800 36118 856
rect 36286 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36670 856
rect 36838 800 36854 856
rect 37022 800 37038 856
rect 37206 800 37222 856
rect 37390 800 37406 856
rect 37574 800 37590 856
rect 37758 800 37774 856
rect 37942 800 37958 856
rect 38126 800 38142 856
rect 38310 800 38326 856
rect 38494 800 38510 856
rect 38678 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39062 856
rect 39230 800 39246 856
rect 39414 800 39430 856
rect 39598 800 39614 856
rect 39782 800 39798 856
rect 39966 800 39982 856
rect 40150 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40534 856
rect 40702 800 40718 856
rect 40886 800 40902 856
rect 41070 800 41086 856
rect 41254 800 41270 856
rect 41438 800 41454 856
rect 41622 800 41638 856
rect 41806 800 41822 856
rect 41990 800 42006 856
rect 42174 800 42190 856
rect 42358 800 42374 856
rect 42542 800 42558 856
rect 42726 800 42742 856
rect 42910 800 42926 856
rect 43094 800 43110 856
rect 43278 800 43294 856
rect 43462 800 43478 856
rect 43646 800 43662 856
rect 43830 800 43846 856
rect 44014 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44398 856
rect 44566 800 44582 856
rect 44750 800 44766 856
rect 44934 800 44950 856
rect 45118 800 45134 856
rect 45302 800 45318 856
rect 45486 800 45502 856
rect 45670 800 45686 856
rect 45854 800 45870 856
rect 46038 800 46054 856
rect 46222 800 46238 856
rect 46406 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46790 856
rect 46958 800 46974 856
rect 47142 800 47158 856
rect 47326 800 47342 856
rect 47510 800 47526 856
rect 47694 800 47710 856
rect 47878 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48262 856
rect 48430 800 48446 856
rect 48614 800 48630 856
rect 48798 800 48814 856
rect 48982 800 48998 856
rect 49166 800 49182 856
rect 49350 800 49366 856
rect 49534 800 49550 856
rect 49718 800 49734 856
rect 49902 800 49918 856
rect 50086 800 50102 856
rect 50270 800 50286 856
rect 50454 800 50470 856
rect 50638 800 50654 856
rect 50822 800 50838 856
rect 51006 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51390 856
rect 51558 800 51574 856
rect 51742 800 51758 856
rect 51926 800 51942 856
rect 52110 800 52126 856
rect 52294 800 52310 856
rect 52478 800 52494 856
rect 52662 800 52678 856
rect 52846 800 52862 856
rect 53030 800 53046 856
rect 53214 800 53230 856
rect 53398 800 53414 856
rect 53582 800 53598 856
rect 53766 800 53782 856
rect 53950 800 53966 856
rect 54134 800 54150 856
rect 54318 800 54334 856
rect 54502 800 54518 856
rect 54686 800 54702 856
rect 54870 800 54886 856
rect 55054 800 55070 856
rect 55238 800 55254 856
rect 55422 800 55438 856
rect 55606 800 55622 856
rect 55790 800 55806 856
rect 55974 800 55990 856
rect 56158 800 56174 856
rect 56342 800 56358 856
rect 56526 800 56542 856
rect 56710 800 56726 856
rect 56894 800 56910 856
rect 57078 800 57094 856
rect 57262 800 57278 856
rect 57446 800 57462 856
rect 57630 800 57646 856
rect 57814 800 57830 856
rect 57998 800 58014 856
rect 58182 800 58198 856
rect 58366 800 58382 856
rect 58550 800 58566 856
rect 58734 800 58750 856
rect 58918 800 58934 856
rect 59102 800 59118 856
rect 59286 800 59302 856
rect 59470 800 59486 856
rect 59654 800 59670 856
rect 59838 800 59854 856
rect 60022 800 60038 856
rect 60206 800 60222 856
rect 60390 800 60406 856
rect 60574 800 60590 856
rect 60758 800 60774 856
rect 60942 800 60958 856
rect 61126 800 61142 856
rect 61310 800 61326 856
rect 61494 800 61510 856
rect 61678 800 61694 856
rect 61862 800 61878 856
rect 62046 800 62062 856
rect 62230 800 62246 856
rect 62414 800 62430 856
rect 62598 800 62614 856
rect 62782 800 62798 856
rect 62966 800 62982 856
rect 63150 800 63166 856
rect 63334 800 63350 856
rect 63518 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63902 856
rect 64070 800 64086 856
rect 64254 800 64270 856
rect 64438 800 64454 856
rect 64622 800 64638 856
rect 64806 800 64822 856
rect 64990 800 65006 856
rect 65174 800 65190 856
rect 65358 800 65374 856
rect 65542 800 65558 856
rect 65726 800 65742 856
rect 65910 800 65926 856
rect 66094 800 66110 856
rect 66278 800 66294 856
rect 66462 800 66478 856
rect 66646 800 66662 856
rect 66830 800 66846 856
rect 67014 800 67030 856
rect 67198 800 67214 856
rect 67382 800 67398 856
rect 67566 800 67582 856
rect 67750 800 67766 856
rect 67934 800 67950 856
rect 68118 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68502 856
rect 68670 800 68686 856
rect 68854 800 68870 856
rect 69038 800 69054 856
rect 69222 800 69238 856
rect 69406 800 69422 856
rect 69590 800 69606 856
rect 69774 800 69790 856
rect 69958 800 69974 856
rect 70142 800 70158 856
rect 70326 800 70342 856
rect 70510 800 70526 856
rect 70694 800 70710 856
rect 70878 800 70894 856
rect 71062 800 71078 856
rect 71246 800 71262 856
rect 71430 800 71446 856
rect 71614 800 71630 856
rect 71798 800 71814 856
rect 71982 800 71998 856
rect 72166 800 72182 856
rect 72350 800 72366 856
rect 72534 800 72550 856
rect 72718 800 72734 856
rect 72902 800 72918 856
rect 73086 800 73102 856
rect 73270 800 73286 856
rect 73454 800 73470 856
rect 73638 800 73654 856
rect 73822 800 73838 856
rect 74006 800 74022 856
rect 74190 800 74206 856
rect 74374 800 74390 856
rect 74558 800 74574 856
rect 74742 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75126 856
rect 75294 800 75310 856
rect 75478 800 75494 856
rect 75662 800 75678 856
rect 75846 800 75862 856
rect 76030 800 76046 856
rect 76214 800 76230 856
rect 76398 800 76414 856
rect 76582 800 76598 856
rect 76766 800 76782 856
rect 76950 800 76966 856
rect 77134 800 77150 856
rect 77318 800 77334 856
rect 77502 800 77518 856
rect 77686 800 77702 856
rect 77870 800 77886 856
rect 78054 800 78070 856
rect 78238 800 78254 856
rect 78422 800 78438 856
rect 78606 800 78622 856
rect 78790 800 78806 856
rect 78974 800 78990 856
rect 79158 800 79174 856
rect 79342 800 79358 856
rect 79526 800 79542 856
rect 79710 800 79726 856
rect 79894 800 79910 856
rect 80078 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80646 856
rect 80814 800 80830 856
rect 80998 800 81014 856
rect 81182 800 81198 856
rect 81366 800 81382 856
rect 81550 800 81566 856
rect 81734 800 81750 856
rect 81918 800 81934 856
rect 82102 800 82118 856
rect 82286 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82670 856
rect 82838 800 82854 856
rect 83022 800 83038 856
rect 83206 800 83222 856
rect 83390 800 83406 856
rect 83574 800 83590 856
rect 83758 800 83774 856
rect 83942 800 83958 856
rect 84126 800 84142 856
rect 84310 800 84326 856
rect 84494 800 84510 856
rect 84678 800 84694 856
rect 84862 800 84878 856
rect 85046 800 85062 856
rect 85230 800 85246 856
rect 85414 800 85430 856
rect 85598 800 85614 856
rect 85782 800 85798 856
rect 85966 800 85982 856
rect 86150 800 86166 856
rect 86334 800 86350 856
rect 86518 800 86534 856
rect 86702 800 86718 856
rect 86886 800 86902 856
rect 87070 800 87086 856
rect 87254 800 87270 856
rect 87438 800 87454 856
rect 87622 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88006 856
rect 88174 800 88190 856
rect 88358 800 88374 856
rect 88542 800 88558 856
rect 88726 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89110 856
rect 89278 800 89294 856
rect 89462 800 89478 856
rect 89646 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90030 856
rect 90198 800 90214 856
rect 90382 800 90398 856
rect 90566 800 90582 856
rect 90750 800 90766 856
rect 90934 800 90950 856
rect 91118 800 91134 856
rect 91302 800 91318 856
rect 91486 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91870 856
rect 92038 800 92054 856
rect 92222 800 92238 856
rect 92406 800 92422 856
rect 92590 800 92606 856
rect 92774 800 92790 856
rect 92958 800 92974 856
rect 93142 800 93158 856
rect 93326 800 93342 856
rect 93510 800 93526 856
rect 93694 800 93710 856
rect 93878 800 93894 856
rect 94062 800 94078 856
rect 94246 800 94262 856
rect 94430 800 94446 856
rect 94614 800 94630 856
rect 94798 800 94814 856
rect 94982 800 94998 856
rect 95166 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95734 856
rect 95902 800 95918 856
rect 96086 800 96102 856
rect 96270 800 96286 856
rect 96454 800 96470 856
rect 96638 800 96654 856
rect 96822 800 96838 856
rect 97006 800 97022 856
rect 97190 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97758 856
rect 97926 800 97942 856
rect 98110 800 98126 856
rect 98294 800 98310 856
rect 98478 800 98494 856
rect 98662 800 98678 856
rect 98846 800 98862 856
rect 99030 800 99046 856
rect 99214 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
rect 99950 800 99966 856
rect 100134 800 100150 856
rect 100318 800 100334 856
rect 100502 800 100518 856
rect 100686 800 100702 856
rect 100870 800 100886 856
rect 101054 800 101070 856
rect 101238 800 101254 856
rect 101422 800 101438 856
rect 101606 800 101622 856
rect 101790 800 101806 856
rect 101974 800 101990 856
rect 102158 800 102174 856
rect 102342 800 102358 856
rect 102526 800 102542 856
rect 102710 800 102726 856
rect 102894 800 102910 856
rect 103078 800 103094 856
rect 103262 800 103278 856
rect 103446 800 103462 856
rect 103630 800 103646 856
rect 103814 800 103830 856
rect 103998 800 104014 856
rect 104182 800 104198 856
rect 104366 800 104382 856
rect 104550 800 104566 856
rect 104734 800 104750 856
rect 104918 800 104934 856
rect 105102 800 105118 856
rect 105286 800 117742 856
<< metal3 >>
rect 0 157904 800 158024
rect 119200 157632 120000 157752
rect 0 154096 800 154216
rect 119200 154096 120000 154216
rect 119200 150560 120000 150680
rect 0 150288 800 150408
rect 119200 147024 120000 147144
rect 0 146480 800 146600
rect 119200 143488 120000 143608
rect 0 142672 800 142792
rect 119200 139952 120000 140072
rect 0 138864 800 138984
rect 119200 136416 120000 136536
rect 0 135056 800 135176
rect 119200 132880 120000 133000
rect 0 131248 800 131368
rect 119200 129344 120000 129464
rect 0 127440 800 127560
rect 119200 125808 120000 125928
rect 0 123632 800 123752
rect 119200 122272 120000 122392
rect 0 119824 800 119944
rect 119200 118736 120000 118856
rect 0 116016 800 116136
rect 119200 115200 120000 115320
rect 0 112208 800 112328
rect 119200 111664 120000 111784
rect 0 108400 800 108520
rect 119200 108128 120000 108248
rect 0 104592 800 104712
rect 119200 104592 120000 104712
rect 119200 101056 120000 101176
rect 0 100784 800 100904
rect 119200 97520 120000 97640
rect 0 96976 800 97096
rect 119200 93984 120000 94104
rect 0 93168 800 93288
rect 119200 90448 120000 90568
rect 0 89360 800 89480
rect 119200 86912 120000 87032
rect 0 85552 800 85672
rect 119200 83376 120000 83496
rect 0 81744 800 81864
rect 119200 79840 120000 79960
rect 0 77936 800 78056
rect 119200 76304 120000 76424
rect 0 74128 800 74248
rect 119200 72768 120000 72888
rect 0 70320 800 70440
rect 119200 69232 120000 69352
rect 0 66512 800 66632
rect 119200 65696 120000 65816
rect 0 62704 800 62824
rect 119200 62160 120000 62280
rect 0 58896 800 59016
rect 119200 58624 120000 58744
rect 0 55088 800 55208
rect 119200 55088 120000 55208
rect 119200 51552 120000 51672
rect 0 51280 800 51400
rect 119200 48016 120000 48136
rect 0 47472 800 47592
rect 119200 44480 120000 44600
rect 0 43664 800 43784
rect 119200 40944 120000 41064
rect 0 39856 800 39976
rect 119200 37408 120000 37528
rect 0 36048 800 36168
rect 119200 33872 120000 33992
rect 0 32240 800 32360
rect 119200 30336 120000 30456
rect 0 28432 800 28552
rect 119200 26800 120000 26920
rect 0 24624 800 24744
rect 119200 23264 120000 23384
rect 0 20816 800 20936
rect 119200 19728 120000 19848
rect 0 17008 800 17128
rect 119200 16192 120000 16312
rect 0 13200 800 13320
rect 119200 12656 120000 12776
rect 0 9392 800 9512
rect 119200 9120 120000 9240
rect 0 5584 800 5704
rect 119200 5584 120000 5704
rect 119200 2048 120000 2168
rect 0 1776 800 1896
<< obsm3 >>
rect 800 157552 119120 157793
rect 800 154296 119200 157552
rect 880 154016 119120 154296
rect 800 150760 119200 154016
rect 800 150488 119120 150760
rect 880 150480 119120 150488
rect 880 150208 119200 150480
rect 800 147224 119200 150208
rect 800 146944 119120 147224
rect 800 146680 119200 146944
rect 880 146400 119200 146680
rect 800 143688 119200 146400
rect 800 143408 119120 143688
rect 800 142872 119200 143408
rect 880 142592 119200 142872
rect 800 140152 119200 142592
rect 800 139872 119120 140152
rect 800 139064 119200 139872
rect 880 138784 119200 139064
rect 800 136616 119200 138784
rect 800 136336 119120 136616
rect 800 135256 119200 136336
rect 880 134976 119200 135256
rect 800 133080 119200 134976
rect 800 132800 119120 133080
rect 800 131448 119200 132800
rect 880 131168 119200 131448
rect 800 129544 119200 131168
rect 800 129264 119120 129544
rect 800 127640 119200 129264
rect 880 127360 119200 127640
rect 800 126008 119200 127360
rect 800 125728 119120 126008
rect 800 123832 119200 125728
rect 880 123552 119200 123832
rect 800 122472 119200 123552
rect 800 122192 119120 122472
rect 800 120024 119200 122192
rect 880 119744 119200 120024
rect 800 118936 119200 119744
rect 800 118656 119120 118936
rect 800 116216 119200 118656
rect 880 115936 119200 116216
rect 800 115400 119200 115936
rect 800 115120 119120 115400
rect 800 112408 119200 115120
rect 880 112128 119200 112408
rect 800 111864 119200 112128
rect 800 111584 119120 111864
rect 800 108600 119200 111584
rect 880 108328 119200 108600
rect 880 108320 119120 108328
rect 800 108048 119120 108320
rect 800 104792 119200 108048
rect 880 104512 119120 104792
rect 800 101256 119200 104512
rect 800 100984 119120 101256
rect 880 100976 119120 100984
rect 880 100704 119200 100976
rect 800 97720 119200 100704
rect 800 97440 119120 97720
rect 800 97176 119200 97440
rect 880 96896 119200 97176
rect 800 94184 119200 96896
rect 800 93904 119120 94184
rect 800 93368 119200 93904
rect 880 93088 119200 93368
rect 800 90648 119200 93088
rect 800 90368 119120 90648
rect 800 89560 119200 90368
rect 880 89280 119200 89560
rect 800 87112 119200 89280
rect 800 86832 119120 87112
rect 800 85752 119200 86832
rect 880 85472 119200 85752
rect 800 83576 119200 85472
rect 800 83296 119120 83576
rect 800 81944 119200 83296
rect 880 81664 119200 81944
rect 800 80040 119200 81664
rect 800 79760 119120 80040
rect 800 78136 119200 79760
rect 880 77856 119200 78136
rect 800 76504 119200 77856
rect 800 76224 119120 76504
rect 800 74328 119200 76224
rect 880 74048 119200 74328
rect 800 72968 119200 74048
rect 800 72688 119120 72968
rect 800 70520 119200 72688
rect 880 70240 119200 70520
rect 800 69432 119200 70240
rect 800 69152 119120 69432
rect 800 66712 119200 69152
rect 880 66432 119200 66712
rect 800 65896 119200 66432
rect 800 65616 119120 65896
rect 800 62904 119200 65616
rect 880 62624 119200 62904
rect 800 62360 119200 62624
rect 800 62080 119120 62360
rect 800 59096 119200 62080
rect 880 58824 119200 59096
rect 880 58816 119120 58824
rect 800 58544 119120 58816
rect 800 55288 119200 58544
rect 880 55008 119120 55288
rect 800 51752 119200 55008
rect 800 51480 119120 51752
rect 880 51472 119120 51480
rect 880 51200 119200 51472
rect 800 48216 119200 51200
rect 800 47936 119120 48216
rect 800 47672 119200 47936
rect 880 47392 119200 47672
rect 800 44680 119200 47392
rect 800 44400 119120 44680
rect 800 43864 119200 44400
rect 880 43584 119200 43864
rect 800 41144 119200 43584
rect 800 40864 119120 41144
rect 800 40056 119200 40864
rect 880 39776 119200 40056
rect 800 37608 119200 39776
rect 800 37328 119120 37608
rect 800 36248 119200 37328
rect 880 35968 119200 36248
rect 800 34072 119200 35968
rect 800 33792 119120 34072
rect 800 32440 119200 33792
rect 880 32160 119200 32440
rect 800 30536 119200 32160
rect 800 30256 119120 30536
rect 800 28632 119200 30256
rect 880 28352 119200 28632
rect 800 27000 119200 28352
rect 800 26720 119120 27000
rect 800 24824 119200 26720
rect 880 24544 119200 24824
rect 800 23464 119200 24544
rect 800 23184 119120 23464
rect 800 21016 119200 23184
rect 880 20736 119200 21016
rect 800 19928 119200 20736
rect 800 19648 119120 19928
rect 800 17208 119200 19648
rect 880 16928 119200 17208
rect 800 16392 119200 16928
rect 800 16112 119120 16392
rect 800 13400 119200 16112
rect 880 13120 119200 13400
rect 800 12856 119200 13120
rect 800 12576 119120 12856
rect 800 9592 119200 12576
rect 880 9320 119200 9592
rect 880 9312 119120 9320
rect 800 9040 119120 9312
rect 800 5784 119200 9040
rect 880 5504 119120 5784
rect 800 2248 119200 5504
rect 800 1976 119120 2248
rect 880 1968 119120 1976
rect 880 1803 119200 1968
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
<< labels >>
rlabel metal3 s 119200 2048 120000 2168 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 119200 108128 120000 108248 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 119200 118736 120000 118856 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 119200 129344 120000 129464 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 119200 139952 120000 140072 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 119200 150560 120000 150680 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 117318 159200 117374 160000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 104070 159200 104126 160000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 90822 159200 90878 160000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 77574 159200 77630 160000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 64326 159200 64382 160000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 119200 12656 120000 12776 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 51078 159200 51134 160000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 37830 159200 37886 160000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 24582 159200 24638 160000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 11334 159200 11390 160000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 157904 800 158024 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 146480 800 146600 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 123632 800 123752 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 100784 800 100904 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 119200 23264 120000 23384 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 89360 800 89480 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 66512 800 66632 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 119200 33872 120000 33992 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 119200 44480 120000 44600 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 119200 55088 120000 55208 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 119200 65696 120000 65816 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 119200 76304 120000 76424 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 119200 86912 120000 87032 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 119200 97520 120000 97640 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 119200 9120 120000 9240 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 119200 115200 120000 115320 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 119200 125808 120000 125928 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 119200 136416 120000 136536 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 119200 147024 120000 147144 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 119200 157632 120000 157752 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 108486 159200 108542 160000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 95238 159200 95294 160000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 81990 159200 82046 160000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 68742 159200 68798 160000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 55494 159200 55550 160000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 119200 19728 120000 19848 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 42246 159200 42302 160000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 28998 159200 29054 160000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 15750 159200 15806 160000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 2502 159200 2558 160000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 150288 800 150408 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 138864 800 138984 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 127440 800 127560 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 116016 800 116136 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 104592 800 104712 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 119200 30336 120000 30456 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 81744 800 81864 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 58896 800 59016 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 47472 800 47592 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 119200 40944 120000 41064 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 119200 51552 120000 51672 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 119200 62160 120000 62280 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 119200 72768 120000 72888 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 119200 83376 120000 83496 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 119200 93984 120000 94104 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 119200 104592 120000 104712 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 119200 5584 120000 5704 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 119200 111664 120000 111784 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 119200 122272 120000 122392 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 119200 132880 120000 133000 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 119200 143488 120000 143608 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 119200 154096 120000 154216 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 112902 159200 112958 160000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 99654 159200 99710 160000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 86406 159200 86462 160000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 73158 159200 73214 160000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 59910 159200 59966 160000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 119200 16192 120000 16312 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 46662 159200 46718 160000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 33414 159200 33470 160000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 20166 159200 20222 160000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 6918 159200 6974 160000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 154096 800 154216 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 142672 800 142792 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 119824 800 119944 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 119200 26800 120000 26920 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 85552 800 85672 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 62704 800 62824 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 119200 37408 120000 37528 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 119200 48016 120000 48136 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 119200 58624 120000 58744 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 119200 69232 120000 69352 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 119200 79840 120000 79960 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 119200 90448 120000 90568 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 119200 101056 120000 101176 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 105174 0 105230 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 14646 0 14702 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6587314
string GDS_FILE /home/kaya/Desktop/caravel_example/caravel_example/openlane/user_proj_example/runs/22_12_02_05_33/results/signoff/user_proj_example.magic.gds
string GDS_START 138062
<< end >>

