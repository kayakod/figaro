magic
tech sky130A
magscale 1 2
timestamp 1659698180
<< metal1 >>
rect 88334 702992 88340 703044
rect 88392 703032 88398 703044
rect 89530 703032 89536 703044
rect 88392 703004 89536 703032
rect 88392 702992 88398 703004
rect 89530 702992 89536 703004
rect 89588 702992 89594 703044
rect 309134 700884 309140 700936
rect 309192 700924 309198 700936
rect 364794 700924 364800 700936
rect 309192 700896 364800 700924
rect 309192 700884 309198 700896
rect 364794 700884 364800 700896
rect 364852 700884 364858 700936
rect 313274 700816 313280 700868
rect 313332 700856 313338 700868
rect 397178 700856 397184 700868
rect 313332 700828 397184 700856
rect 313332 700816 313338 700828
rect 397178 700816 397184 700828
rect 397236 700816 397242 700868
rect 317414 700748 317420 700800
rect 317472 700788 317478 700800
rect 413370 700788 413376 700800
rect 317472 700760 413376 700788
rect 317472 700748 317478 700760
rect 413370 700748 413376 700760
rect 413428 700748 413434 700800
rect 321554 700680 321560 700732
rect 321612 700720 321618 700732
rect 429562 700720 429568 700732
rect 321612 700692 429568 700720
rect 321612 700680 321618 700692
rect 429562 700680 429568 700692
rect 429620 700680 429626 700732
rect 327074 700612 327080 700664
rect 327132 700652 327138 700664
rect 461946 700652 461952 700664
rect 327132 700624 461952 700652
rect 327132 700612 327138 700624
rect 461946 700612 461952 700624
rect 462004 700612 462010 700664
rect 331306 700544 331312 700596
rect 331364 700584 331370 700596
rect 478138 700584 478144 700596
rect 331364 700556 478144 700584
rect 331364 700544 331370 700556
rect 478138 700544 478144 700556
rect 478196 700544 478202 700596
rect 295334 700476 295340 700528
rect 295392 700516 295398 700528
rect 300026 700516 300032 700528
rect 295392 700488 300032 700516
rect 295392 700476 295398 700488
rect 300026 700476 300032 700488
rect 300084 700476 300090 700528
rect 335354 700476 335360 700528
rect 335412 700516 335418 700528
rect 494330 700516 494336 700528
rect 335412 700488 494336 700516
rect 335412 700476 335418 700488
rect 494330 700476 494336 700488
rect 494388 700476 494394 700528
rect 339494 700408 339500 700460
rect 339552 700448 339558 700460
rect 526714 700448 526720 700460
rect 339552 700420 526720 700448
rect 339552 700408 339558 700420
rect 526714 700408 526720 700420
rect 526772 700408 526778 700460
rect 299474 700340 299480 700392
rect 299532 700380 299538 700392
rect 332410 700380 332416 700392
rect 299532 700352 332416 700380
rect 299532 700340 299538 700352
rect 332410 700340 332416 700352
rect 332468 700340 332474 700392
rect 343634 700340 343640 700392
rect 343692 700380 343698 700392
rect 542906 700380 542912 700392
rect 343692 700352 542912 700380
rect 343692 700340 343698 700352
rect 542906 700340 542912 700352
rect 542964 700340 542970 700392
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 279418 700312 279424 700324
rect 267700 700284 279424 700312
rect 267700 700272 267706 700284
rect 279418 700272 279424 700284
rect 279476 700272 279482 700324
rect 304994 700272 305000 700324
rect 305052 700312 305058 700324
rect 348602 700312 348608 700324
rect 305052 700284 348608 700312
rect 305052 700272 305058 700284
rect 348602 700272 348608 700284
rect 348660 700272 348666 700324
rect 349154 700272 349160 700324
rect 349212 700312 349218 700324
rect 559098 700312 559104 700324
rect 349212 700284 559104 700312
rect 349212 700272 349218 700284
rect 559098 700272 559104 700284
rect 559156 700272 559162 700324
rect 23474 697552 23480 697604
rect 23532 697592 23538 697604
rect 24762 697592 24768 697604
rect 23532 697564 24768 697592
rect 23532 697552 23538 697564
rect 24762 697552 24768 697564
rect 24820 697552 24826 697604
rect 2774 680552 2780 680604
rect 2832 680592 2838 680604
rect 4798 680592 4804 680604
rect 2832 680564 4804 680592
rect 2832 680552 2838 680564
rect 4798 680552 4804 680564
rect 4856 680552 4862 680604
rect 353938 680348 353944 680400
rect 353996 680388 354002 680400
rect 580166 680388 580172 680400
rect 353996 680360 580172 680388
rect 353996 680348 354002 680360
rect 580166 680348 580172 680360
rect 580224 680348 580230 680400
rect 360838 667904 360844 667956
rect 360896 667944 360902 667956
rect 580166 667944 580172 667956
rect 360896 667916 580172 667944
rect 360896 667904 360902 667916
rect 580166 667904 580172 667916
rect 580224 667904 580230 667956
rect 367738 641724 367744 641776
rect 367796 641764 367802 641776
rect 579890 641764 579896 641776
rect 367796 641736 579896 641764
rect 367796 641724 367802 641736
rect 579890 641724 579896 641736
rect 579948 641724 579954 641776
rect 3602 629280 3608 629332
rect 3660 629320 3666 629332
rect 35158 629320 35164 629332
rect 3660 629292 35164 629320
rect 3660 629280 3666 629292
rect 35158 629280 35164 629292
rect 35216 629280 35222 629332
rect 377398 627920 377404 627972
rect 377456 627960 377462 627972
rect 579890 627960 579896 627972
rect 377456 627932 579896 627960
rect 377456 627920 377462 627932
rect 579890 627920 579896 627932
rect 579948 627920 579954 627972
rect 3326 615476 3332 615528
rect 3384 615516 3390 615528
rect 22738 615516 22744 615528
rect 3384 615488 22744 615516
rect 3384 615476 3390 615488
rect 22738 615476 22744 615488
rect 22796 615476 22802 615528
rect 509878 615476 509884 615528
rect 509936 615516 509942 615528
rect 580166 615516 580172 615528
rect 509936 615488 580172 615516
rect 509936 615476 509942 615488
rect 580166 615476 580172 615488
rect 580224 615476 580230 615528
rect 3326 603100 3332 603152
rect 3384 603140 3390 603152
rect 14458 603140 14464 603152
rect 3384 603112 14464 603140
rect 3384 603100 3390 603112
rect 14458 603100 14464 603112
rect 14516 603100 14522 603152
rect 3326 576852 3332 576904
rect 3384 576892 3390 576904
rect 7558 576892 7564 576904
rect 3384 576864 7564 576892
rect 3384 576852 3390 576864
rect 7558 576852 7564 576864
rect 7616 576852 7622 576904
rect 359458 561688 359464 561740
rect 359516 561728 359522 561740
rect 580166 561728 580172 561740
rect 359516 561700 580172 561728
rect 359516 561688 359522 561700
rect 580166 561688 580172 561700
rect 580224 561688 580230 561740
rect 364978 535440 364984 535492
rect 365036 535480 365042 535492
rect 580166 535480 580172 535492
rect 365036 535452 580172 535480
rect 365036 535440 365042 535452
rect 580166 535440 580172 535452
rect 580224 535440 580230 535492
rect 3326 525784 3332 525836
rect 3384 525824 3390 525836
rect 61378 525824 61384 525836
rect 3384 525796 61384 525824
rect 3384 525784 3390 525796
rect 61378 525784 61384 525796
rect 61436 525784 61442 525836
rect 374638 522996 374644 523048
rect 374696 523036 374702 523048
rect 580166 523036 580172 523048
rect 374696 523008 580172 523036
rect 374696 522996 374702 523008
rect 580166 522996 580172 523008
rect 580224 522996 580230 523048
rect 3326 513340 3332 513392
rect 3384 513380 3390 513392
rect 25498 513380 25504 513392
rect 3384 513352 25504 513380
rect 3384 513340 3390 513352
rect 25498 513340 25504 513352
rect 25556 513340 25562 513392
rect 356698 509260 356704 509312
rect 356756 509300 356762 509312
rect 579614 509300 579620 509312
rect 356756 509272 579620 509300
rect 356756 509260 356762 509272
rect 579614 509260 579620 509272
rect 579672 509260 579678 509312
rect 2958 499536 2964 499588
rect 3016 499576 3022 499588
rect 17218 499576 17224 499588
rect 3016 499548 17224 499576
rect 3016 499536 3022 499548
rect 17218 499536 17224 499548
rect 17276 499536 17282 499588
rect 3234 474036 3240 474088
rect 3292 474076 3298 474088
rect 8938 474076 8944 474088
rect 3292 474048 8944 474076
rect 3292 474036 3298 474048
rect 8938 474036 8944 474048
rect 8996 474036 9002 474088
rect 355318 456764 355324 456816
rect 355376 456804 355382 456816
rect 580166 456804 580172 456816
rect 355376 456776 580172 456804
rect 355376 456764 355382 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 373258 430584 373264 430636
rect 373316 430624 373322 430636
rect 579798 430624 579804 430636
rect 373316 430596 579804 430624
rect 373316 430584 373322 430596
rect 579798 430584 579804 430596
rect 579856 430584 579862 430636
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 180058 422328 180064 422340
rect 3016 422300 180064 422328
rect 3016 422288 3022 422300
rect 180058 422288 180064 422300
rect 180116 422288 180122 422340
rect 381538 416780 381544 416832
rect 381596 416820 381602 416832
rect 579614 416820 579620 416832
rect 381596 416792 579620 416820
rect 381596 416780 381602 416792
rect 579614 416780 579620 416792
rect 579672 416780 579678 416832
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 26878 409884 26884 409896
rect 3384 409856 26884 409884
rect 3384 409844 3390 409856
rect 26878 409844 26884 409856
rect 26936 409844 26942 409896
rect 363598 404336 363604 404388
rect 363656 404376 363662 404388
rect 580166 404376 580172 404388
rect 363656 404348 580172 404376
rect 363656 404336 363662 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 2958 396040 2964 396092
rect 3016 396080 3022 396092
rect 18598 396080 18604 396092
rect 3016 396052 18604 396080
rect 3016 396040 3022 396052
rect 18598 396040 18604 396052
rect 18656 396040 18662 396092
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 10318 371260 10324 371272
rect 3384 371232 10324 371260
rect 3384 371220 3390 371232
rect 10318 371220 10324 371232
rect 10376 371220 10382 371272
rect 354030 364352 354036 364404
rect 354088 364392 354094 364404
rect 580166 364392 580172 364404
rect 354088 364364 580172 364392
rect 354088 364352 354094 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 371878 324300 371884 324352
rect 371936 324340 371942 324352
rect 580166 324340 580172 324352
rect 371936 324312 580172 324340
rect 371936 324300 371942 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 224218 318832 224224 318844
rect 3384 318804 224224 318832
rect 3384 318792 3390 318804
rect 224218 318792 224224 318804
rect 224276 318792 224282 318844
rect 378778 311856 378784 311908
rect 378836 311896 378842 311908
rect 580166 311896 580172 311908
rect 378836 311868 580172 311896
rect 378836 311856 378842 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3326 306348 3332 306400
rect 3384 306388 3390 306400
rect 28258 306388 28264 306400
rect 3384 306360 28264 306388
rect 3384 306348 3390 306360
rect 28258 306348 28264 306360
rect 28316 306348 28322 306400
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 21358 292584 21364 292596
rect 3384 292556 21364 292584
rect 3384 292544 3390 292556
rect 21358 292544 21364 292556
rect 21416 292544 21422 292596
rect 369118 271872 369124 271924
rect 369176 271912 369182 271924
rect 579982 271912 579988 271924
rect 369176 271884 579988 271912
rect 369176 271872 369182 271884
rect 579982 271872 579988 271884
rect 580040 271872 580046 271924
rect 3326 267724 3332 267776
rect 3384 267764 3390 267776
rect 13078 267764 13084 267776
rect 3384 267736 13084 267764
rect 3384 267724 3390 267736
rect 13078 267724 13084 267736
rect 13136 267724 13142 267776
rect 218054 263508 218060 263560
rect 218112 263548 218118 263560
rect 278682 263548 278688 263560
rect 218112 263520 278688 263548
rect 218112 263508 218118 263520
rect 278682 263508 278688 263520
rect 278740 263508 278746 263560
rect 202874 263440 202880 263492
rect 202932 263480 202938 263492
rect 274266 263480 274272 263492
rect 202932 263452 274272 263480
rect 202932 263440 202938 263452
rect 274266 263440 274272 263452
rect 274324 263440 274330 263492
rect 169754 263372 169760 263424
rect 169812 263412 169818 263424
rect 269850 263412 269856 263424
rect 169812 263384 269856 263412
rect 169812 263372 169818 263384
rect 269850 263372 269856 263384
rect 269908 263372 269914 263424
rect 153194 263304 153200 263356
rect 153252 263344 153258 263356
rect 265434 263344 265440 263356
rect 153252 263316 265440 263344
rect 153252 263304 153258 263316
rect 265434 263304 265440 263316
rect 265492 263304 265498 263356
rect 138014 263236 138020 263288
rect 138072 263276 138078 263288
rect 261018 263276 261024 263288
rect 138072 263248 261024 263276
rect 138072 263236 138078 263248
rect 261018 263236 261024 263248
rect 261076 263236 261082 263288
rect 104894 263168 104900 263220
rect 104952 263208 104958 263220
rect 256602 263208 256608 263220
rect 104952 263180 256608 263208
rect 104952 263168 104958 263180
rect 256602 263168 256608 263180
rect 256660 263168 256666 263220
rect 88334 263100 88340 263152
rect 88392 263140 88398 263152
rect 252186 263140 252192 263152
rect 88392 263112 252192 263140
rect 88392 263100 88398 263112
rect 252186 263100 252192 263112
rect 252244 263100 252250 263152
rect 73154 263032 73160 263084
rect 73212 263072 73218 263084
rect 247770 263072 247776 263084
rect 73212 263044 247776 263072
rect 73212 263032 73218 263044
rect 247770 263032 247776 263044
rect 247828 263032 247834 263084
rect 40034 262964 40040 263016
rect 40092 263004 40098 263016
rect 243354 263004 243360 263016
rect 40092 262976 243360 263004
rect 40092 262964 40098 262976
rect 243354 262964 243360 262976
rect 243412 262964 243418 263016
rect 282914 262964 282920 263016
rect 282972 263004 282978 263016
rect 291930 263004 291936 263016
rect 282972 262976 291936 263004
rect 282972 262964 282978 262976
rect 291930 262964 291936 262976
rect 291988 262964 291994 263016
rect 23474 262896 23480 262948
rect 23532 262936 23538 262948
rect 238938 262936 238944 262948
rect 23532 262908 238944 262936
rect 23532 262896 23538 262908
rect 238938 262896 238944 262908
rect 238996 262896 239002 262948
rect 279418 262896 279424 262948
rect 279476 262936 279482 262948
rect 287514 262936 287520 262948
rect 279476 262908 287520 262936
rect 279476 262896 279482 262908
rect 287514 262896 287520 262908
rect 287572 262896 287578 262948
rect 8294 262828 8300 262880
rect 8352 262868 8358 262880
rect 234522 262868 234528 262880
rect 8352 262840 234528 262868
rect 8352 262828 8358 262840
rect 234522 262828 234528 262840
rect 234580 262828 234586 262880
rect 234614 262828 234620 262880
rect 234672 262868 234678 262880
rect 283098 262868 283104 262880
rect 234672 262840 283104 262868
rect 234672 262828 234678 262840
rect 283098 262828 283104 262840
rect 283156 262828 283162 262880
rect 354122 259428 354128 259480
rect 354180 259468 354186 259480
rect 580166 259468 580172 259480
rect 354180 259440 580172 259468
rect 354180 259428 354186 259440
rect 580166 259428 580172 259440
rect 580224 259428 580230 259480
rect 4798 258000 4804 258052
rect 4856 258040 4862 258052
rect 230382 258040 230388 258052
rect 4856 258012 230388 258040
rect 4856 258000 4862 258012
rect 230382 258000 230388 258012
rect 230440 258000 230446 258052
rect 353294 258000 353300 258052
rect 353352 258040 353358 258052
rect 580166 258040 580172 258052
rect 353352 258012 580172 258040
rect 353352 258000 353358 258012
rect 580166 258000 580172 258012
rect 580224 258000 580230 258052
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 230382 255252 230388 255264
rect 3476 255224 230388 255252
rect 3476 255212 3482 255224
rect 230382 255212 230388 255224
rect 230440 255212 230446 255264
rect 3510 251132 3516 251184
rect 3568 251172 3574 251184
rect 230382 251172 230388 251184
rect 3568 251144 230388 251172
rect 3568 251132 3574 251144
rect 230382 251132 230388 251144
rect 230440 251132 230446 251184
rect 353294 251132 353300 251184
rect 353352 251172 353358 251184
rect 360838 251172 360844 251184
rect 353352 251144 360844 251172
rect 353352 251132 353358 251144
rect 360838 251132 360844 251144
rect 360896 251132 360902 251184
rect 353294 248344 353300 248396
rect 353352 248384 353358 248396
rect 367738 248384 367744 248396
rect 353352 248356 367744 248384
rect 353352 248344 353358 248356
rect 367738 248344 367744 248356
rect 367796 248344 367802 248396
rect 35158 246984 35164 247036
rect 35216 247024 35222 247036
rect 229646 247024 229652 247036
rect 35216 246996 229652 247024
rect 35216 246984 35222 246996
rect 229646 246984 229652 246996
rect 229704 246984 229710 247036
rect 353294 244196 353300 244248
rect 353352 244236 353358 244248
rect 377398 244236 377404 244248
rect 353352 244208 377404 244236
rect 353352 244196 353358 244208
rect 377398 244196 377404 244208
rect 377456 244196 377462 244248
rect 22738 242836 22744 242888
rect 22796 242876 22802 242888
rect 229278 242876 229284 242888
rect 22796 242848 229284 242876
rect 22796 242836 22802 242848
rect 229278 242836 229284 242848
rect 229336 242836 229342 242888
rect 14458 240048 14464 240100
rect 14516 240088 14522 240100
rect 230014 240088 230020 240100
rect 14516 240060 230020 240088
rect 14516 240048 14522 240060
rect 230014 240048 230020 240060
rect 230072 240048 230078 240100
rect 353294 240048 353300 240100
rect 353352 240088 353358 240100
rect 509878 240088 509884 240100
rect 353352 240060 509884 240088
rect 353352 240048 353358 240060
rect 509878 240048 509884 240060
rect 509936 240048 509942 240100
rect 353294 237328 353300 237380
rect 353352 237368 353358 237380
rect 580350 237368 580356 237380
rect 353352 237340 580356 237368
rect 353352 237328 353358 237340
rect 580350 237328 580356 237340
rect 580408 237328 580414 237380
rect 7558 235900 7564 235952
rect 7616 235940 7622 235952
rect 230198 235940 230204 235952
rect 7616 235912 230204 235940
rect 7616 235900 7622 235912
rect 230198 235900 230204 235912
rect 230256 235900 230262 235952
rect 353294 233180 353300 233232
rect 353352 233220 353358 233232
rect 580442 233220 580448 233232
rect 353352 233192 580448 233220
rect 353352 233180 353358 233192
rect 580442 233180 580448 233192
rect 580500 233180 580506 233232
rect 3602 231752 3608 231804
rect 3660 231792 3666 231804
rect 230382 231792 230388 231804
rect 3660 231764 230388 231792
rect 3660 231752 3666 231764
rect 230382 231752 230388 231764
rect 230440 231752 230446 231804
rect 353294 230392 353300 230444
rect 353352 230432 353358 230444
rect 359458 230432 359464 230444
rect 353352 230404 359464 230432
rect 353352 230392 353358 230404
rect 359458 230392 359464 230404
rect 359516 230392 359522 230444
rect 3694 227672 3700 227724
rect 3752 227712 3758 227724
rect 230382 227712 230388 227724
rect 3752 227684 230388 227712
rect 3752 227672 3758 227684
rect 230382 227672 230388 227684
rect 230440 227672 230446 227724
rect 353294 226244 353300 226296
rect 353352 226284 353358 226296
rect 364978 226284 364984 226296
rect 353352 226256 364984 226284
rect 353352 226244 353358 226256
rect 364978 226244 364984 226256
rect 365036 226244 365042 226296
rect 61378 224884 61384 224936
rect 61436 224924 61442 224936
rect 229646 224924 229652 224936
rect 61436 224896 229652 224924
rect 61436 224884 61442 224896
rect 229646 224884 229652 224896
rect 229704 224884 229710 224936
rect 353294 223524 353300 223576
rect 353352 223564 353358 223576
rect 374638 223564 374644 223576
rect 353352 223536 374644 223564
rect 353352 223524 353358 223536
rect 374638 223524 374644 223536
rect 374696 223524 374702 223576
rect 25498 220736 25504 220788
rect 25556 220776 25562 220788
rect 230382 220776 230388 220788
rect 25556 220748 230388 220776
rect 25556 220736 25562 220748
rect 230382 220736 230388 220748
rect 230440 220736 230446 220788
rect 353938 219444 353944 219496
rect 353996 219484 354002 219496
rect 580166 219484 580172 219496
rect 353996 219456 580172 219484
rect 353996 219444 354002 219456
rect 580166 219444 580172 219456
rect 580224 219444 580230 219496
rect 353294 219376 353300 219428
rect 353352 219416 353358 219428
rect 356698 219416 356704 219428
rect 353352 219388 356704 219416
rect 353352 219376 353358 219388
rect 356698 219376 356704 219388
rect 356756 219376 356762 219428
rect 17218 216588 17224 216640
rect 17276 216628 17282 216640
rect 230382 216628 230388 216640
rect 17276 216600 230388 216628
rect 17276 216588 17282 216600
rect 230382 216588 230388 216600
rect 230440 216588 230446 216640
rect 353294 215228 353300 215280
rect 353352 215268 353358 215280
rect 580534 215268 580540 215280
rect 353352 215240 580540 215268
rect 353352 215228 353358 215240
rect 580534 215228 580540 215240
rect 580592 215228 580598 215280
rect 8938 212440 8944 212492
rect 8996 212480 9002 212492
rect 230382 212480 230388 212492
rect 8996 212452 230388 212480
rect 8996 212440 9002 212452
rect 230382 212440 230388 212452
rect 230440 212440 230446 212492
rect 353294 212440 353300 212492
rect 353352 212480 353358 212492
rect 580626 212480 580632 212492
rect 353352 212452 580632 212480
rect 353352 212440 353358 212452
rect 580626 212440 580632 212452
rect 580684 212440 580690 212492
rect 3786 209720 3792 209772
rect 3844 209760 3850 209772
rect 229646 209760 229652 209772
rect 3844 209732 229652 209760
rect 3844 209720 3850 209732
rect 229646 209720 229652 209732
rect 229704 209720 229710 209772
rect 353294 208156 353300 208208
rect 353352 208196 353358 208208
rect 355318 208196 355324 208208
rect 353352 208168 355324 208196
rect 353352 208156 353358 208168
rect 355318 208156 355324 208168
rect 355376 208156 355382 208208
rect 3878 205572 3884 205624
rect 3936 205612 3942 205624
rect 229462 205612 229468 205624
rect 3936 205584 229468 205612
rect 3936 205572 3942 205584
rect 229462 205572 229468 205584
rect 229520 205572 229526 205624
rect 353294 205572 353300 205624
rect 353352 205612 353358 205624
rect 373258 205612 373264 205624
rect 353352 205584 373264 205612
rect 353352 205572 353358 205584
rect 373258 205572 373264 205584
rect 373316 205572 373322 205624
rect 180058 201424 180064 201476
rect 180116 201464 180122 201476
rect 230382 201464 230388 201476
rect 180116 201436 230388 201464
rect 180116 201424 180122 201436
rect 230382 201424 230388 201436
rect 230440 201424 230446 201476
rect 353294 201424 353300 201476
rect 353352 201464 353358 201476
rect 381538 201464 381544 201476
rect 353352 201436 381544 201464
rect 353352 201424 353358 201436
rect 381538 201424 381544 201436
rect 381596 201424 381602 201476
rect 353294 198636 353300 198688
rect 353352 198676 353358 198688
rect 363598 198676 363604 198688
rect 353352 198648 363604 198676
rect 353352 198636 353358 198648
rect 363598 198636 363604 198648
rect 363656 198636 363662 198688
rect 26878 197276 26884 197328
rect 26936 197316 26942 197328
rect 229830 197316 229836 197328
rect 26936 197288 229836 197316
rect 26936 197276 26942 197288
rect 229830 197276 229836 197288
rect 229888 197276 229894 197328
rect 353294 194488 353300 194540
rect 353352 194528 353358 194540
rect 580718 194528 580724 194540
rect 353352 194500 580724 194528
rect 353352 194488 353358 194500
rect 580718 194488 580724 194500
rect 580776 194488 580782 194540
rect 18598 193128 18604 193180
rect 18656 193168 18662 193180
rect 230382 193168 230388 193180
rect 18656 193140 230388 193168
rect 18656 193128 18662 193140
rect 230382 193128 230388 193140
rect 230440 193128 230446 193180
rect 10318 190408 10324 190460
rect 10376 190448 10382 190460
rect 230382 190448 230388 190460
rect 10376 190420 230388 190448
rect 10376 190408 10382 190420
rect 230382 190408 230388 190420
rect 230440 190408 230446 190460
rect 353294 187620 353300 187672
rect 353352 187660 353358 187672
rect 580810 187660 580816 187672
rect 353352 187632 580816 187660
rect 353352 187620 353358 187632
rect 580810 187620 580816 187632
rect 580868 187620 580874 187672
rect 3970 186260 3976 186312
rect 4028 186300 4034 186312
rect 230382 186300 230388 186312
rect 4028 186272 230388 186300
rect 4028 186260 4034 186272
rect 230382 186260 230388 186272
rect 230440 186260 230446 186312
rect 353294 183472 353300 183524
rect 353352 183512 353358 183524
rect 371878 183512 371884 183524
rect 353352 183484 371884 183512
rect 353352 183472 353358 183484
rect 371878 183472 371884 183484
rect 371936 183472 371942 183524
rect 4062 182112 4068 182164
rect 4120 182152 4126 182164
rect 229830 182152 229836 182164
rect 4120 182124 229836 182152
rect 4120 182112 4126 182124
rect 229830 182112 229836 182124
rect 229888 182112 229894 182164
rect 353294 180752 353300 180804
rect 353352 180792 353358 180804
rect 378778 180792 378784 180804
rect 353352 180764 378784 180792
rect 353352 180752 353358 180764
rect 378778 180752 378784 180764
rect 378836 180752 378842 180804
rect 354030 179392 354036 179444
rect 354088 179432 354094 179444
rect 579614 179432 579620 179444
rect 354088 179404 579620 179432
rect 354088 179392 354094 179404
rect 579614 179392 579620 179404
rect 579672 179392 579678 179444
rect 224218 177964 224224 178016
rect 224276 178004 224282 178016
rect 230382 178004 230388 178016
rect 224276 177976 230388 178004
rect 224276 177964 224282 177976
rect 230382 177964 230388 177976
rect 230440 177964 230446 178016
rect 353294 176604 353300 176656
rect 353352 176644 353358 176656
rect 580902 176644 580908 176656
rect 353352 176616 580908 176644
rect 353352 176604 353358 176616
rect 580902 176604 580908 176616
rect 580960 176604 580966 176656
rect 28258 175176 28264 175228
rect 28316 175216 28322 175228
rect 230382 175216 230388 175228
rect 28316 175188 230388 175216
rect 28316 175176 28322 175188
rect 230382 175176 230388 175188
rect 230440 175176 230446 175228
rect 353294 173816 353300 173868
rect 353352 173856 353358 173868
rect 369118 173856 369124 173868
rect 353352 173828 369124 173856
rect 353352 173816 353358 173828
rect 369118 173816 369124 173828
rect 369176 173816 369182 173868
rect 21358 171028 21364 171080
rect 21416 171068 21422 171080
rect 230382 171068 230388 171080
rect 21416 171040 230388 171068
rect 21416 171028 21422 171040
rect 230382 171028 230388 171040
rect 230440 171028 230446 171080
rect 13078 166948 13084 167000
rect 13136 166988 13142 167000
rect 230382 166988 230388 167000
rect 13136 166960 230388 166988
rect 13136 166948 13142 166960
rect 230382 166948 230388 166960
rect 230440 166948 230446 167000
rect 353294 166948 353300 167000
rect 353352 166988 353358 167000
rect 580258 166988 580264 167000
rect 353352 166960 580264 166988
rect 353352 166948 353358 166960
rect 580258 166948 580264 166960
rect 580316 166948 580322 167000
rect 3326 162800 3332 162852
rect 3384 162840 3390 162852
rect 230382 162840 230388 162852
rect 3384 162812 230388 162840
rect 3384 162800 3390 162812
rect 230382 162800 230388 162812
rect 230440 162800 230446 162852
rect 353294 162800 353300 162852
rect 353352 162840 353358 162852
rect 580350 162840 580356 162852
rect 353352 162812 580356 162840
rect 353352 162800 353358 162812
rect 580350 162800 580356 162812
rect 580408 162800 580414 162852
rect 3418 160012 3424 160064
rect 3476 160052 3482 160064
rect 230382 160052 230388 160064
rect 3476 160024 230388 160052
rect 3476 160012 3482 160024
rect 230382 160012 230388 160024
rect 230440 160012 230446 160064
rect 3510 155864 3516 155916
rect 3568 155904 3574 155916
rect 229278 155904 229284 155916
rect 3568 155876 229284 155904
rect 3568 155864 3574 155876
rect 229278 155864 229284 155876
rect 229336 155864 229342 155916
rect 353294 155864 353300 155916
rect 353352 155904 353358 155916
rect 580442 155904 580448 155916
rect 353352 155876 580448 155904
rect 353352 155864 353358 155876
rect 580442 155864 580448 155876
rect 580500 155864 580506 155916
rect 353938 153212 353944 153264
rect 353996 153252 354002 153264
rect 579614 153252 579620 153264
rect 353996 153224 579620 153252
rect 353996 153212 354002 153224
rect 579614 153212 579620 153224
rect 579672 153212 579678 153264
rect 3602 151716 3608 151768
rect 3660 151756 3666 151768
rect 230382 151756 230388 151768
rect 3660 151728 230388 151756
rect 3660 151716 3666 151728
rect 230382 151716 230388 151728
rect 230440 151716 230446 151768
rect 353294 151716 353300 151768
rect 353352 151756 353358 151768
rect 580534 151756 580540 151768
rect 353352 151728 580540 151756
rect 353352 151716 353358 151728
rect 580534 151716 580540 151728
rect 580592 151716 580598 151768
rect 3694 147568 3700 147620
rect 3752 147608 3758 147620
rect 230382 147608 230388 147620
rect 3752 147580 230388 147608
rect 3752 147568 3758 147580
rect 230382 147568 230388 147580
rect 230440 147568 230446 147620
rect 3786 144848 3792 144900
rect 3844 144888 3850 144900
rect 230014 144888 230020 144900
rect 3844 144860 230020 144888
rect 3844 144848 3850 144860
rect 230014 144848 230020 144860
rect 230072 144848 230078 144900
rect 353294 144848 353300 144900
rect 353352 144888 353358 144900
rect 580626 144888 580632 144900
rect 353352 144860 580632 144888
rect 353352 144848 353358 144860
rect 580626 144848 580632 144860
rect 580684 144848 580690 144900
rect 353294 140768 353300 140820
rect 353352 140808 353358 140820
rect 580166 140808 580172 140820
rect 353352 140780 580172 140808
rect 353352 140768 353358 140780
rect 580166 140768 580172 140780
rect 580224 140768 580230 140820
rect 3418 140700 3424 140752
rect 3476 140740 3482 140752
rect 230382 140740 230388 140752
rect 3476 140712 230388 140740
rect 3476 140700 3482 140712
rect 230382 140700 230388 140712
rect 230440 140700 230446 140752
rect 3418 136552 3424 136604
rect 3476 136592 3482 136604
rect 229646 136592 229652 136604
rect 3476 136564 229652 136592
rect 3476 136552 3482 136564
rect 229646 136552 229652 136564
rect 229704 136552 229710 136604
rect 3602 128324 3608 128376
rect 3660 128364 3666 128376
rect 230382 128364 230388 128376
rect 3660 128336 230388 128364
rect 3660 128324 3666 128336
rect 230382 128324 230388 128336
rect 230440 128324 230446 128376
rect 354214 128256 354220 128308
rect 354272 128296 354278 128308
rect 580166 128296 580172 128308
rect 354272 128268 580172 128296
rect 354272 128256 354278 128268
rect 580166 128256 580172 128268
rect 580224 128256 580230 128308
rect 3510 115948 3516 116000
rect 3568 115988 3574 116000
rect 230382 115988 230388 116000
rect 3568 115960 230388 115988
rect 3568 115948 3574 115960
rect 230382 115948 230388 115960
rect 230440 115948 230446 116000
rect 353938 114452 353944 114504
rect 353996 114492 354002 114504
rect 580166 114492 580172 114504
rect 353996 114464 580172 114492
rect 353996 114452 354002 114464
rect 580166 114452 580172 114464
rect 580224 114452 580230 114504
rect 3142 113092 3148 113144
rect 3200 113132 3206 113144
rect 229738 113132 229744 113144
rect 3200 113104 229744 113132
rect 3200 113092 3206 113104
rect 229738 113092 229744 113104
rect 229796 113092 229802 113144
rect 3418 104864 3424 104916
rect 3476 104904 3482 104916
rect 230382 104904 230388 104916
rect 3476 104876 230388 104904
rect 3476 104864 3482 104876
rect 230382 104864 230388 104876
rect 230440 104864 230446 104916
rect 354582 102076 354588 102128
rect 354640 102116 354646 102128
rect 579982 102116 579988 102128
rect 354640 102088 579988 102116
rect 354640 102076 354646 102088
rect 579982 102076 579988 102088
rect 580040 102076 580046 102128
rect 247678 97928 247684 97980
rect 247736 97968 247742 97980
rect 248506 97968 248512 97980
rect 247736 97940 248512 97968
rect 247736 97928 247742 97940
rect 248506 97928 248512 97940
rect 248564 97928 248570 97980
rect 286318 97928 286324 97980
rect 286376 97968 286382 97980
rect 287330 97968 287336 97980
rect 286376 97940 287336 97968
rect 286376 97928 286382 97940
rect 287330 97928 287336 97940
rect 287388 97928 287394 97980
rect 303890 97928 303896 97980
rect 303948 97968 303954 97980
rect 307110 97968 307116 97980
rect 303948 97940 307116 97968
rect 303948 97928 303954 97940
rect 307110 97928 307116 97940
rect 307168 97928 307174 97980
rect 246942 97860 246948 97912
rect 247000 97900 247006 97912
rect 249978 97900 249984 97912
rect 247000 97872 249984 97900
rect 247000 97860 247006 97872
rect 249978 97860 249984 97872
rect 250036 97860 250042 97912
rect 276750 97860 276756 97912
rect 276808 97900 276814 97912
rect 277762 97900 277768 97912
rect 276808 97872 277768 97900
rect 276808 97860 276814 97872
rect 277762 97860 277768 97872
rect 277820 97860 277826 97912
rect 284938 97860 284944 97912
rect 284996 97900 285002 97912
rect 287146 97900 287152 97912
rect 284996 97872 287152 97900
rect 284996 97860 285002 97872
rect 287146 97860 287152 97872
rect 287204 97860 287210 97912
rect 332962 97860 332968 97912
rect 333020 97900 333026 97912
rect 338758 97900 338764 97912
rect 333020 97872 338764 97900
rect 333020 97860 333026 97872
rect 338758 97860 338764 97872
rect 338816 97860 338822 97912
rect 244918 97792 244924 97844
rect 244976 97832 244982 97844
rect 255682 97832 255688 97844
rect 244976 97804 255688 97832
rect 244976 97792 244982 97804
rect 255682 97792 255688 97804
rect 255740 97792 255746 97844
rect 282270 97792 282276 97844
rect 282328 97832 282334 97844
rect 288802 97832 288808 97844
rect 282328 97804 288808 97832
rect 282328 97792 282334 97804
rect 288802 97792 288808 97804
rect 288860 97792 288866 97844
rect 294138 97792 294144 97844
rect 294196 97832 294202 97844
rect 300302 97832 300308 97844
rect 294196 97804 300308 97832
rect 294196 97792 294202 97804
rect 300302 97792 300308 97804
rect 300360 97792 300366 97844
rect 334618 97792 334624 97844
rect 334676 97832 334682 97844
rect 337470 97832 337476 97844
rect 334676 97804 337476 97832
rect 334676 97792 334682 97804
rect 337470 97792 337476 97804
rect 337528 97792 337534 97844
rect 235258 97724 235264 97776
rect 235316 97764 235322 97776
rect 249242 97764 249248 97776
rect 235316 97736 249248 97764
rect 235316 97724 235322 97736
rect 249242 97724 249248 97736
rect 249300 97724 249306 97776
rect 294874 97724 294880 97776
rect 294932 97764 294938 97776
rect 301774 97764 301780 97776
rect 294932 97736 301780 97764
rect 294932 97724 294938 97736
rect 301774 97724 301780 97736
rect 301832 97724 301838 97776
rect 325786 97724 325792 97776
rect 325844 97764 325850 97776
rect 339034 97764 339040 97776
rect 325844 97736 339040 97764
rect 325844 97724 325850 97736
rect 339034 97724 339040 97736
rect 339092 97724 339098 97776
rect 243538 97656 243544 97708
rect 243596 97696 243602 97708
rect 266170 97696 266176 97708
rect 243596 97668 266176 97696
rect 243596 97656 243602 97668
rect 266170 97656 266176 97668
rect 266228 97656 266234 97708
rect 293954 97656 293960 97708
rect 294012 97696 294018 97708
rect 300854 97696 300860 97708
rect 294012 97668 300860 97696
rect 294012 97656 294018 97668
rect 300854 97656 300860 97668
rect 300912 97656 300918 97708
rect 316402 97656 316408 97708
rect 316460 97696 316466 97708
rect 326338 97696 326344 97708
rect 316460 97668 326344 97696
rect 316460 97656 316466 97668
rect 326338 97656 326344 97668
rect 326396 97656 326402 97708
rect 330754 97656 330760 97708
rect 330812 97696 330818 97708
rect 347038 97696 347044 97708
rect 330812 97668 347044 97696
rect 330812 97656 330818 97668
rect 347038 97656 347044 97668
rect 347096 97656 347102 97708
rect 242158 97588 242164 97640
rect 242216 97628 242222 97640
rect 272242 97628 272248 97640
rect 242216 97600 272248 97628
rect 242216 97588 242222 97600
rect 272242 97588 272248 97600
rect 272300 97588 272306 97640
rect 278406 97588 278412 97640
rect 278464 97628 278470 97640
rect 281074 97628 281080 97640
rect 278464 97600 281080 97628
rect 278464 97588 278470 97600
rect 281074 97588 281080 97600
rect 281132 97588 281138 97640
rect 295610 97588 295616 97640
rect 295668 97628 295674 97640
rect 304534 97628 304540 97640
rect 295668 97600 304540 97628
rect 295668 97588 295674 97600
rect 304534 97588 304540 97600
rect 304592 97588 304598 97640
rect 321922 97588 321928 97640
rect 321980 97628 321986 97640
rect 338850 97628 338856 97640
rect 321980 97600 338856 97628
rect 321980 97588 321986 97600
rect 338850 97588 338856 97600
rect 338908 97588 338914 97640
rect 239398 97520 239404 97572
rect 239456 97560 239462 97572
rect 274450 97560 274456 97572
rect 239456 97532 274456 97560
rect 239456 97520 239462 97532
rect 274450 97520 274456 97532
rect 274508 97520 274514 97572
rect 279878 97520 279884 97572
rect 279936 97560 279942 97572
rect 289354 97560 289360 97572
rect 279936 97532 289360 97560
rect 279936 97520 279942 97532
rect 289354 97520 289360 97532
rect 289412 97520 289418 97572
rect 294322 97520 294328 97572
rect 294380 97560 294386 97572
rect 303614 97560 303620 97572
rect 294380 97532 303620 97560
rect 294380 97520 294386 97532
rect 303614 97520 303620 97532
rect 303672 97520 303678 97572
rect 322474 97520 322480 97572
rect 322532 97560 322538 97572
rect 341518 97560 341524 97572
rect 322532 97532 341524 97560
rect 322532 97520 322538 97532
rect 341518 97520 341524 97532
rect 341576 97520 341582 97572
rect 128354 97452 128360 97504
rect 128412 97492 128418 97504
rect 264882 97492 264888 97504
rect 128412 97464 264888 97492
rect 128412 97452 128418 97464
rect 264882 97452 264888 97464
rect 264940 97452 264946 97504
rect 275278 97452 275284 97504
rect 275336 97492 275342 97504
rect 285674 97492 285680 97504
rect 275336 97464 285680 97492
rect 275336 97452 275342 97464
rect 285674 97452 285680 97464
rect 285732 97452 285738 97504
rect 299290 97452 299296 97504
rect 299348 97492 299354 97504
rect 322934 97492 322940 97504
rect 299348 97464 322940 97492
rect 299348 97452 299354 97464
rect 322934 97452 322940 97464
rect 322992 97452 322998 97504
rect 324682 97452 324688 97504
rect 324740 97492 324746 97504
rect 342898 97492 342904 97504
rect 324740 97464 342904 97492
rect 324740 97452 324746 97464
rect 342898 97452 342904 97464
rect 342956 97452 342962 97504
rect 238018 97384 238024 97436
rect 238076 97424 238082 97436
rect 281626 97424 281632 97436
rect 238076 97396 281632 97424
rect 238076 97384 238082 97396
rect 281626 97384 281632 97396
rect 281684 97384 281690 97436
rect 288434 97424 288440 97436
rect 287026 97396 288440 97424
rect 121454 97316 121460 97368
rect 121512 97356 121518 97368
rect 263778 97356 263784 97368
rect 121512 97328 263784 97356
rect 121512 97316 121518 97328
rect 263778 97316 263784 97328
rect 263836 97316 263842 97368
rect 278038 97316 278044 97368
rect 278096 97356 278102 97368
rect 287026 97356 287054 97396
rect 288434 97384 288440 97396
rect 288492 97384 288498 97436
rect 298186 97384 298192 97436
rect 298244 97424 298250 97436
rect 324038 97424 324044 97436
rect 298244 97396 324044 97424
rect 298244 97384 298250 97396
rect 324038 97384 324044 97396
rect 324096 97384 324102 97436
rect 326890 97384 326896 97436
rect 326948 97424 326954 97436
rect 345658 97424 345664 97436
rect 326948 97396 345664 97424
rect 326948 97384 326954 97396
rect 345658 97384 345664 97396
rect 345716 97384 345722 97436
rect 278096 97328 287054 97356
rect 278096 97316 278102 97328
rect 297082 97316 297088 97368
rect 297140 97356 297146 97368
rect 320910 97356 320916 97368
rect 297140 97328 320916 97356
rect 297140 97316 297146 97328
rect 320910 97316 320916 97328
rect 320968 97316 320974 97368
rect 321370 97316 321376 97368
rect 321428 97356 321434 97368
rect 349798 97356 349804 97368
rect 321428 97328 349804 97356
rect 321428 97316 321434 97328
rect 349798 97316 349804 97328
rect 349856 97316 349862 97368
rect 28258 97248 28264 97300
rect 28316 97288 28322 97300
rect 247586 97288 247592 97300
rect 28316 97260 247592 97288
rect 28316 97248 28322 97260
rect 247586 97248 247592 97260
rect 247644 97248 247650 97300
rect 273990 97248 273996 97300
rect 274048 97288 274054 97300
rect 274048 97260 277394 97288
rect 274048 97248 274054 97260
rect 264974 97180 264980 97232
rect 265032 97220 265038 97232
rect 272794 97220 272800 97232
rect 265032 97192 272800 97220
rect 265032 97180 265038 97192
rect 272794 97180 272800 97192
rect 272852 97180 272858 97232
rect 277366 97220 277394 97260
rect 278222 97248 278228 97300
rect 278280 97288 278286 97300
rect 279050 97288 279056 97300
rect 278280 97260 279056 97288
rect 278280 97248 278286 97260
rect 279050 97248 279056 97260
rect 279108 97248 279114 97300
rect 286042 97288 286048 97300
rect 281460 97260 286048 97288
rect 281460 97220 281488 97260
rect 286042 97248 286048 97260
rect 286100 97248 286106 97300
rect 297634 97248 297640 97300
rect 297692 97288 297698 97300
rect 323486 97288 323492 97300
rect 297692 97260 323492 97288
rect 297692 97248 297698 97260
rect 323486 97248 323492 97260
rect 323544 97248 323550 97300
rect 326430 97248 326436 97300
rect 326488 97288 326494 97300
rect 475378 97288 475384 97300
rect 326488 97260 475384 97288
rect 326488 97248 326494 97260
rect 475378 97248 475384 97260
rect 475436 97248 475442 97300
rect 277366 97192 281488 97220
rect 281534 97180 281540 97232
rect 281592 97220 281598 97232
rect 283282 97220 283288 97232
rect 281592 97192 283288 97220
rect 281592 97180 281598 97192
rect 283282 97180 283288 97192
rect 283340 97180 283346 97232
rect 330202 97180 330208 97232
rect 330260 97220 330266 97232
rect 338942 97220 338948 97232
rect 330260 97192 338948 97220
rect 330260 97180 330266 97192
rect 338942 97180 338948 97192
rect 339000 97180 339006 97232
rect 255958 97112 255964 97164
rect 256016 97152 256022 97164
rect 258442 97152 258448 97164
rect 256016 97124 258448 97152
rect 256016 97112 256022 97124
rect 258442 97112 258448 97124
rect 258500 97112 258506 97164
rect 257430 96976 257436 97028
rect 257488 97016 257494 97028
rect 258994 97016 259000 97028
rect 257488 96988 259000 97016
rect 257488 96976 257494 96988
rect 258994 96976 259000 96988
rect 259052 96976 259058 97028
rect 261018 96976 261024 97028
rect 261076 97016 261082 97028
rect 261478 97016 261484 97028
rect 261076 96988 261484 97016
rect 261076 96976 261082 96988
rect 261478 96976 261484 96988
rect 261536 96976 261542 97028
rect 274174 96976 274180 97028
rect 274232 97016 274238 97028
rect 277210 97016 277216 97028
rect 274232 96988 277216 97016
rect 274232 96976 274238 96988
rect 277210 96976 277216 96988
rect 277268 96976 277274 97028
rect 265158 96908 265164 96960
rect 265216 96948 265222 96960
rect 265618 96948 265624 96960
rect 265216 96920 265624 96948
rect 265216 96908 265222 96920
rect 265618 96908 265624 96920
rect 265676 96908 265682 96960
rect 273622 96908 273628 96960
rect 273680 96948 273686 96960
rect 274082 96948 274088 96960
rect 273680 96920 274088 96948
rect 273680 96908 273686 96920
rect 274082 96908 274088 96920
rect 274140 96908 274146 96960
rect 275094 96908 275100 96960
rect 275152 96948 275158 96960
rect 275370 96948 275376 96960
rect 275152 96920 275376 96948
rect 275152 96908 275158 96920
rect 275370 96908 275376 96920
rect 275428 96908 275434 96960
rect 279602 96908 279608 96960
rect 279660 96948 279666 96960
rect 280522 96948 280528 96960
rect 279660 96920 280528 96948
rect 279660 96908 279666 96920
rect 280522 96908 280528 96920
rect 280580 96908 280586 96960
rect 287146 96908 287152 96960
rect 287204 96948 287210 96960
rect 287698 96948 287704 96960
rect 287204 96920 287704 96948
rect 287204 96908 287210 96920
rect 287698 96908 287704 96920
rect 287756 96908 287762 96960
rect 289170 96908 289176 96960
rect 289228 96948 289234 96960
rect 289906 96948 289912 96960
rect 289228 96920 289912 96948
rect 289228 96908 289234 96920
rect 289906 96908 289912 96920
rect 289964 96908 289970 96960
rect 335722 96908 335728 96960
rect 335780 96948 335786 96960
rect 337378 96948 337384 96960
rect 335780 96920 337384 96948
rect 335780 96908 335786 96920
rect 337378 96908 337384 96920
rect 337436 96908 337442 96960
rect 243630 96840 243636 96892
rect 243688 96880 243694 96892
rect 247034 96880 247040 96892
rect 243688 96852 247040 96880
rect 243688 96840 243694 96852
rect 247034 96840 247040 96852
rect 247092 96840 247098 96892
rect 264238 96840 264244 96892
rect 264296 96880 264302 96892
rect 266722 96880 266728 96892
rect 264296 96852 266728 96880
rect 264296 96840 264302 96852
rect 266722 96840 266728 96852
rect 266780 96840 266786 96892
rect 272518 96840 272524 96892
rect 272576 96880 272582 96892
rect 274818 96880 274824 96892
rect 272576 96852 274824 96880
rect 272576 96840 272582 96852
rect 274818 96840 274824 96852
rect 274876 96840 274882 96892
rect 279694 96840 279700 96892
rect 279752 96880 279758 96892
rect 286594 96880 286600 96892
rect 279752 96852 286600 96880
rect 279752 96840 279758 96852
rect 286594 96840 286600 96852
rect 286652 96840 286658 96892
rect 335354 96840 335360 96892
rect 335412 96880 335418 96892
rect 340138 96880 340144 96892
rect 335412 96852 340144 96880
rect 335412 96840 335418 96852
rect 340138 96840 340144 96852
rect 340196 96840 340202 96892
rect 246390 96772 246396 96824
rect 246448 96812 246454 96824
rect 247770 96812 247776 96824
rect 246448 96784 247776 96812
rect 246448 96772 246454 96784
rect 247770 96772 247776 96784
rect 247828 96772 247834 96824
rect 252922 96772 252928 96824
rect 252980 96812 252986 96824
rect 253106 96812 253112 96824
rect 252980 96784 253112 96812
rect 252980 96772 252986 96784
rect 253106 96772 253112 96784
rect 253164 96772 253170 96824
rect 260926 96772 260932 96824
rect 260984 96812 260990 96824
rect 261386 96812 261392 96824
rect 260984 96784 261392 96812
rect 260984 96772 260990 96784
rect 261386 96772 261392 96784
rect 261444 96772 261450 96824
rect 263686 96772 263692 96824
rect 263744 96812 263750 96824
rect 264146 96812 264152 96824
rect 263744 96784 264152 96812
rect 263744 96772 263750 96784
rect 264146 96772 264152 96784
rect 264204 96772 264210 96824
rect 271138 96772 271144 96824
rect 271196 96812 271202 96824
rect 271874 96812 271880 96824
rect 271196 96784 271880 96812
rect 271196 96772 271202 96784
rect 271874 96772 271880 96784
rect 271932 96772 271938 96824
rect 282178 96772 282184 96824
rect 282236 96812 282242 96824
rect 284846 96812 284852 96824
rect 282236 96784 284852 96812
rect 282236 96772 282242 96784
rect 284846 96772 284852 96784
rect 284904 96772 284910 96824
rect 288618 96772 288624 96824
rect 288676 96812 288682 96824
rect 289078 96812 289084 96824
rect 288676 96784 289084 96812
rect 288676 96772 288682 96784
rect 289078 96772 289084 96784
rect 289136 96772 289142 96824
rect 301130 96772 301136 96824
rect 301188 96812 301194 96824
rect 302970 96812 302976 96824
rect 301188 96784 302976 96812
rect 301188 96772 301194 96784
rect 302970 96772 302976 96784
rect 303028 96772 303034 96824
rect 303614 96772 303620 96824
rect 303672 96812 303678 96824
rect 304258 96812 304264 96824
rect 303672 96784 304264 96812
rect 303672 96772 303678 96784
rect 304258 96772 304264 96784
rect 304316 96772 304322 96824
rect 308122 96772 308128 96824
rect 308180 96812 308186 96824
rect 309778 96812 309784 96824
rect 308180 96784 309784 96812
rect 308180 96772 308186 96784
rect 309778 96772 309784 96784
rect 309836 96772 309842 96824
rect 311986 96772 311992 96824
rect 312044 96812 312050 96824
rect 315298 96812 315304 96824
rect 312044 96784 315304 96812
rect 312044 96772 312050 96784
rect 315298 96772 315304 96784
rect 315356 96772 315362 96824
rect 316954 96772 316960 96824
rect 317012 96812 317018 96824
rect 318058 96812 318064 96824
rect 317012 96784 318064 96812
rect 317012 96772 317018 96784
rect 318058 96772 318064 96784
rect 318116 96772 318122 96824
rect 322934 96772 322940 96824
rect 322992 96812 322998 96824
rect 323762 96812 323768 96824
rect 322992 96784 323768 96812
rect 322992 96772 322998 96784
rect 323762 96772 323768 96784
rect 323820 96772 323826 96824
rect 260098 96704 260104 96756
rect 260156 96744 260162 96756
rect 262306 96744 262312 96756
rect 260156 96716 262312 96744
rect 260156 96704 260162 96716
rect 262306 96704 262312 96716
rect 262364 96704 262370 96756
rect 265618 96704 265624 96756
rect 265676 96744 265682 96756
rect 267274 96744 267280 96756
rect 265676 96716 267280 96744
rect 265676 96704 265682 96716
rect 267274 96704 267280 96716
rect 267332 96704 267338 96756
rect 274082 96704 274088 96756
rect 274140 96744 274146 96756
rect 275002 96744 275008 96756
rect 274140 96716 275008 96744
rect 274140 96704 274146 96716
rect 275002 96704 275008 96716
rect 275060 96704 275066 96756
rect 276658 96704 276664 96756
rect 276716 96744 276722 96756
rect 277578 96744 277584 96756
rect 276716 96716 277584 96744
rect 276716 96704 276722 96716
rect 277578 96704 277584 96716
rect 277636 96704 277642 96756
rect 285858 96744 285864 96756
rect 283576 96716 285864 96744
rect 283576 96688 283604 96716
rect 285858 96704 285864 96716
rect 285916 96704 285922 96756
rect 287698 96704 287704 96756
rect 287756 96744 287762 96756
rect 290458 96744 290464 96756
rect 287756 96716 290464 96744
rect 287756 96704 287762 96716
rect 290458 96704 290464 96716
rect 290516 96704 290522 96756
rect 300854 96704 300860 96756
rect 300912 96744 300918 96756
rect 301498 96744 301504 96756
rect 300912 96716 301504 96744
rect 300912 96704 300918 96716
rect 301498 96704 301504 96716
rect 301556 96704 301562 96756
rect 318794 96704 318800 96756
rect 318852 96744 318858 96756
rect 325050 96744 325056 96756
rect 318852 96716 325056 96744
rect 318852 96704 318858 96716
rect 325050 96704 325056 96716
rect 325108 96704 325114 96756
rect 246298 96636 246304 96688
rect 246356 96676 246362 96688
rect 246942 96676 246948 96688
rect 246356 96648 246948 96676
rect 246356 96636 246362 96648
rect 246942 96636 246948 96648
rect 247000 96636 247006 96688
rect 257338 96636 257344 96688
rect 257396 96676 257402 96688
rect 258074 96676 258080 96688
rect 257396 96648 258080 96676
rect 257396 96636 257402 96648
rect 258074 96636 258080 96648
rect 258132 96636 258138 96688
rect 276106 96676 276112 96688
rect 274652 96648 276112 96676
rect 269390 96568 269396 96620
rect 269448 96608 269454 96620
rect 274652 96608 274680 96648
rect 276106 96636 276112 96648
rect 276164 96636 276170 96688
rect 279418 96636 279424 96688
rect 279476 96676 279482 96688
rect 279878 96676 279884 96688
rect 279476 96648 279884 96676
rect 279476 96636 279482 96648
rect 279878 96636 279884 96648
rect 279936 96636 279942 96688
rect 283098 96636 283104 96688
rect 283156 96676 283162 96688
rect 283466 96676 283472 96688
rect 283156 96648 283472 96676
rect 283156 96636 283162 96648
rect 283466 96636 283472 96648
rect 283524 96636 283530 96688
rect 283558 96636 283564 96688
rect 283616 96636 283622 96688
rect 283650 96636 283656 96688
rect 283708 96676 283714 96688
rect 284570 96676 284576 96688
rect 283708 96648 284576 96676
rect 283708 96636 283714 96648
rect 284570 96636 284576 96648
rect 284628 96636 284634 96688
rect 289078 96636 289084 96688
rect 289136 96676 289142 96688
rect 290090 96676 290096 96688
rect 289136 96648 290096 96676
rect 289136 96636 289142 96648
rect 290090 96636 290096 96648
rect 290148 96636 290154 96688
rect 269448 96580 274680 96608
rect 269448 96568 269454 96580
rect 224954 96228 224960 96280
rect 225012 96268 225018 96280
rect 278406 96268 278412 96280
rect 225012 96240 278412 96268
rect 225012 96228 225018 96240
rect 278406 96228 278412 96240
rect 278464 96228 278470 96280
rect 299842 96228 299848 96280
rect 299900 96268 299906 96280
rect 338114 96268 338120 96280
rect 299900 96240 338120 96268
rect 299900 96228 299906 96240
rect 338114 96228 338120 96240
rect 338172 96228 338178 96280
rect 216674 96160 216680 96212
rect 216732 96200 216738 96212
rect 279510 96200 279516 96212
rect 216732 96172 279516 96200
rect 216732 96160 216738 96172
rect 279510 96160 279516 96172
rect 279568 96160 279574 96212
rect 302602 96160 302608 96212
rect 302660 96200 302666 96212
rect 354674 96200 354680 96212
rect 302660 96172 354680 96200
rect 302660 96160 302666 96172
rect 354674 96160 354680 96172
rect 354732 96160 354738 96212
rect 195974 96092 195980 96144
rect 196032 96132 196038 96144
rect 269390 96132 269396 96144
rect 196032 96104 269396 96132
rect 196032 96092 196038 96104
rect 269390 96092 269396 96104
rect 269448 96092 269454 96144
rect 269482 96092 269488 96144
rect 269540 96132 269546 96144
rect 269666 96132 269672 96144
rect 269540 96104 269672 96132
rect 269540 96092 269546 96104
rect 269666 96092 269672 96104
rect 269724 96092 269730 96144
rect 308674 96092 308680 96144
rect 308732 96132 308738 96144
rect 390554 96132 390560 96144
rect 308732 96104 390560 96132
rect 308732 96092 308738 96104
rect 390554 96092 390560 96104
rect 390612 96092 390618 96144
rect 169754 96024 169760 96076
rect 169812 96064 169818 96076
rect 271690 96064 271696 96076
rect 169812 96036 271696 96064
rect 169812 96024 169818 96036
rect 271690 96024 271696 96036
rect 271748 96024 271754 96076
rect 316034 96024 316040 96076
rect 316092 96064 316098 96076
rect 434714 96064 434720 96076
rect 316092 96036 434720 96064
rect 316092 96024 316098 96036
rect 434714 96024 434720 96036
rect 434772 96024 434778 96076
rect 81434 95956 81440 96008
rect 81492 95996 81498 96008
rect 257154 95996 257160 96008
rect 81492 95968 257160 95996
rect 81492 95956 81498 95968
rect 257154 95956 257160 95968
rect 257212 95956 257218 96008
rect 323026 95956 323032 96008
rect 323084 95996 323090 96008
rect 477494 95996 477500 96008
rect 323084 95968 477500 95996
rect 323084 95956 323090 95968
rect 477494 95956 477500 95968
rect 477552 95956 477558 96008
rect 75914 95888 75920 95940
rect 75972 95928 75978 95940
rect 256234 95928 256240 95940
rect 75972 95900 256240 95928
rect 75972 95888 75978 95900
rect 256234 95888 256240 95900
rect 256292 95888 256298 95940
rect 327442 95888 327448 95940
rect 327500 95928 327506 95940
rect 503714 95928 503720 95940
rect 327500 95900 503720 95928
rect 327500 95888 327506 95900
rect 503714 95888 503720 95900
rect 503772 95888 503778 95940
rect 277854 95684 277860 95736
rect 277912 95724 277918 95736
rect 278130 95724 278136 95736
rect 277912 95696 278136 95724
rect 277912 95684 277918 95696
rect 278130 95684 278136 95696
rect 278188 95684 278194 95736
rect 279418 95548 279424 95600
rect 279476 95588 279482 95600
rect 279694 95588 279700 95600
rect 279476 95560 279700 95588
rect 279476 95548 279482 95560
rect 279694 95548 279700 95560
rect 279752 95548 279758 95600
rect 273990 95412 273996 95464
rect 274048 95452 274054 95464
rect 274174 95452 274180 95464
rect 274048 95424 274180 95452
rect 274048 95412 274054 95424
rect 274174 95412 274180 95424
rect 274232 95412 274238 95464
rect 269114 95208 269120 95260
rect 269172 95248 269178 95260
rect 269298 95248 269304 95260
rect 269172 95220 269304 95248
rect 269172 95208 269178 95220
rect 269298 95208 269304 95220
rect 269356 95208 269362 95260
rect 281626 95140 281632 95192
rect 281684 95180 281690 95192
rect 282362 95180 282368 95192
rect 281684 95152 282368 95180
rect 281684 95140 281690 95152
rect 282362 95140 282368 95152
rect 282420 95140 282426 95192
rect 238754 94800 238760 94852
rect 238812 94840 238818 94852
rect 281534 94840 281540 94852
rect 238812 94812 281540 94840
rect 238812 94800 238818 94812
rect 281534 94800 281540 94812
rect 281592 94800 281598 94852
rect 213914 94732 213920 94784
rect 213972 94772 213978 94784
rect 278222 94772 278228 94784
rect 213972 94744 278228 94772
rect 213972 94732 213978 94744
rect 278222 94732 278228 94744
rect 278280 94732 278286 94784
rect 303154 94732 303160 94784
rect 303212 94772 303218 94784
rect 357434 94772 357440 94784
rect 303212 94744 357440 94772
rect 303212 94732 303218 94744
rect 357434 94732 357440 94744
rect 357492 94732 357498 94784
rect 198734 94664 198740 94716
rect 198792 94704 198798 94716
rect 276566 94704 276572 94716
rect 198792 94676 276572 94704
rect 198792 94664 198798 94676
rect 276566 94664 276572 94676
rect 276624 94664 276630 94716
rect 310698 94664 310704 94716
rect 310756 94704 310762 94716
rect 402974 94704 402980 94716
rect 310756 94676 402980 94704
rect 310756 94664 310762 94676
rect 402974 94664 402980 94676
rect 403032 94664 403038 94716
rect 175274 94596 175280 94648
rect 175332 94636 175338 94648
rect 264974 94636 264980 94648
rect 175332 94608 264980 94636
rect 175332 94596 175338 94608
rect 264974 94596 264980 94608
rect 265032 94596 265038 94648
rect 313642 94596 313648 94648
rect 313700 94636 313706 94648
rect 420914 94636 420920 94648
rect 313700 94608 420920 94636
rect 313700 94596 313706 94608
rect 420914 94596 420920 94608
rect 420972 94596 420978 94648
rect 66254 94528 66260 94580
rect 66312 94568 66318 94580
rect 254578 94568 254584 94580
rect 66312 94540 254584 94568
rect 66312 94528 66318 94540
rect 254578 94528 254584 94540
rect 254636 94528 254642 94580
rect 323578 94528 323584 94580
rect 323636 94568 323642 94580
rect 480254 94568 480260 94580
rect 323636 94540 480260 94568
rect 323636 94528 323642 94540
rect 480254 94528 480260 94540
rect 480312 94528 480318 94580
rect 40034 94460 40040 94512
rect 40092 94500 40098 94512
rect 250162 94500 250168 94512
rect 40092 94472 250168 94500
rect 40092 94460 40098 94472
rect 250162 94460 250168 94472
rect 250220 94460 250226 94512
rect 298738 94460 298744 94512
rect 298796 94500 298802 94512
rect 331214 94500 331220 94512
rect 298796 94472 331220 94500
rect 298796 94460 298802 94472
rect 331214 94460 331220 94472
rect 331272 94460 331278 94512
rect 331306 94460 331312 94512
rect 331364 94500 331370 94512
rect 527174 94500 527180 94512
rect 331364 94472 527180 94500
rect 331364 94460 331370 94472
rect 527174 94460 527180 94472
rect 527232 94460 527238 94512
rect 255314 94392 255320 94444
rect 255372 94432 255378 94444
rect 255498 94432 255504 94444
rect 255372 94404 255504 94432
rect 255372 94392 255378 94404
rect 255498 94392 255504 94404
rect 255556 94392 255562 94444
rect 241514 93440 241520 93492
rect 241572 93480 241578 93492
rect 283834 93480 283840 93492
rect 241572 93452 283840 93480
rect 241572 93440 241578 93452
rect 283834 93440 283840 93452
rect 283892 93440 283898 93492
rect 219434 93372 219440 93424
rect 219492 93412 219498 93424
rect 280154 93412 280160 93424
rect 219492 93384 280160 93412
rect 219492 93372 219498 93384
rect 280154 93372 280160 93384
rect 280212 93372 280218 93424
rect 302970 93372 302976 93424
rect 303028 93412 303034 93424
rect 346394 93412 346400 93424
rect 303028 93384 346400 93412
rect 303028 93372 303034 93384
rect 346394 93372 346400 93384
rect 346452 93372 346458 93424
rect 205634 93304 205640 93356
rect 205692 93344 205698 93356
rect 276750 93344 276756 93356
rect 205692 93316 276756 93344
rect 205692 93304 205698 93316
rect 276750 93304 276756 93316
rect 276808 93304 276814 93356
rect 300946 93304 300952 93356
rect 301004 93344 301010 93356
rect 345014 93344 345020 93356
rect 301004 93316 345020 93344
rect 301004 93304 301010 93316
rect 345014 93304 345020 93316
rect 345072 93304 345078 93356
rect 179414 93236 179420 93288
rect 179472 93276 179478 93288
rect 273346 93276 273352 93288
rect 179472 93248 273352 93276
rect 179472 93236 179478 93248
rect 273346 93236 273352 93248
rect 273404 93236 273410 93288
rect 309778 93236 309784 93288
rect 309836 93276 309842 93288
rect 387794 93276 387800 93288
rect 309836 93248 387800 93276
rect 309836 93236 309842 93248
rect 387794 93236 387800 93248
rect 387852 93236 387858 93288
rect 63494 93168 63500 93220
rect 63552 93208 63558 93220
rect 254026 93208 254032 93220
rect 63552 93180 254032 93208
rect 63552 93168 63558 93180
rect 254026 93168 254032 93180
rect 254084 93168 254090 93220
rect 324130 93168 324136 93220
rect 324188 93208 324194 93220
rect 484394 93208 484400 93220
rect 324188 93180 484400 93208
rect 324188 93168 324194 93180
rect 484394 93168 484400 93180
rect 484452 93168 484458 93220
rect 56594 93100 56600 93152
rect 56652 93140 56658 93152
rect 253106 93140 253112 93152
rect 56652 93112 253112 93140
rect 56652 93100 56658 93112
rect 253106 93100 253112 93112
rect 253164 93100 253170 93152
rect 334066 93100 334072 93152
rect 334124 93140 334130 93152
rect 543734 93140 543740 93152
rect 334124 93112 543740 93140
rect 334124 93100 334130 93112
rect 543734 93100 543740 93112
rect 543792 93100 543798 93152
rect 233234 92012 233240 92064
rect 233292 92052 233298 92064
rect 281626 92052 281632 92064
rect 233292 92024 281632 92052
rect 233292 92012 233298 92024
rect 281626 92012 281632 92024
rect 281684 92012 281690 92064
rect 303706 92012 303712 92064
rect 303764 92052 303770 92064
rect 361574 92052 361580 92064
rect 303764 92024 361580 92052
rect 303764 92012 303770 92024
rect 361574 92012 361580 92024
rect 361632 92012 361638 92064
rect 212534 91944 212540 91996
rect 212592 91984 212598 91996
rect 278866 91984 278872 91996
rect 212592 91956 278872 91984
rect 212592 91944 212598 91956
rect 278866 91944 278872 91956
rect 278924 91944 278930 91996
rect 307938 91944 307944 91996
rect 307996 91984 308002 91996
rect 386414 91984 386420 91996
rect 307996 91956 386420 91984
rect 307996 91944 308002 91956
rect 386414 91944 386420 91956
rect 386472 91944 386478 91996
rect 182174 91876 182180 91928
rect 182232 91916 182238 91928
rect 273806 91916 273812 91928
rect 182232 91888 273812 91916
rect 182232 91876 182238 91888
rect 273806 91876 273812 91888
rect 273864 91876 273870 91928
rect 300394 91876 300400 91928
rect 300452 91916 300458 91928
rect 340874 91916 340880 91928
rect 300452 91888 340880 91916
rect 300452 91876 300458 91888
rect 340874 91876 340880 91888
rect 340932 91876 340938 91928
rect 349798 91876 349804 91928
rect 349856 91916 349862 91928
rect 467834 91916 467840 91928
rect 349856 91888 467840 91916
rect 349856 91876 349862 91888
rect 467834 91876 467840 91888
rect 467892 91876 467898 91928
rect 155954 91808 155960 91860
rect 156012 91848 156018 91860
rect 269666 91848 269672 91860
rect 156012 91820 269672 91848
rect 156012 91808 156018 91820
rect 269666 91808 269672 91820
rect 269724 91808 269730 91860
rect 319162 91808 319168 91860
rect 319220 91848 319226 91860
rect 454034 91848 454040 91860
rect 319220 91820 454040 91848
rect 319220 91808 319226 91820
rect 454034 91808 454040 91820
rect 454092 91808 454098 91860
rect 106274 91740 106280 91792
rect 106332 91780 106338 91792
rect 261202 91780 261208 91792
rect 106332 91752 261208 91780
rect 106332 91740 106338 91752
rect 261202 91740 261208 91752
rect 261260 91740 261266 91792
rect 333514 91740 333520 91792
rect 333572 91780 333578 91792
rect 539594 91780 539600 91792
rect 333572 91752 539600 91780
rect 333572 91740 333578 91752
rect 539594 91740 539600 91752
rect 539652 91740 539658 91792
rect 237374 90584 237380 90636
rect 237432 90624 237438 90636
rect 283466 90624 283472 90636
rect 237432 90596 283472 90624
rect 237432 90584 237438 90596
rect 283466 90584 283472 90596
rect 283524 90584 283530 90636
rect 300026 90584 300032 90636
rect 300084 90624 300090 90636
rect 339494 90624 339500 90636
rect 300084 90596 339500 90624
rect 300084 90584 300090 90596
rect 339494 90584 339500 90596
rect 339552 90584 339558 90636
rect 219526 90516 219532 90568
rect 219584 90556 219590 90568
rect 279970 90556 279976 90568
rect 219584 90528 279976 90556
rect 219584 90516 219590 90528
rect 279970 90516 279976 90528
rect 280028 90516 280034 90568
rect 307018 90516 307024 90568
rect 307076 90556 307082 90568
rect 362954 90556 362960 90568
rect 307076 90528 362960 90556
rect 307076 90516 307082 90528
rect 362954 90516 362960 90528
rect 363012 90516 363018 90568
rect 189074 90448 189080 90500
rect 189132 90488 189138 90500
rect 274082 90488 274088 90500
rect 189132 90460 274088 90488
rect 189132 90448 189138 90460
rect 274082 90448 274088 90460
rect 274140 90448 274146 90500
rect 304166 90448 304172 90500
rect 304224 90488 304230 90500
rect 364334 90488 364340 90500
rect 304224 90460 364340 90488
rect 304224 90448 304230 90460
rect 364334 90448 364340 90460
rect 364392 90448 364398 90500
rect 173894 90380 173900 90432
rect 173952 90420 173958 90432
rect 272426 90420 272432 90432
rect 173952 90392 272432 90420
rect 173952 90380 173958 90392
rect 272426 90380 272432 90392
rect 272484 90380 272490 90432
rect 325234 90380 325240 90432
rect 325292 90420 325298 90432
rect 489914 90420 489920 90432
rect 325292 90392 489920 90420
rect 325292 90380 325298 90392
rect 489914 90380 489920 90392
rect 489972 90380 489978 90432
rect 92474 90312 92480 90364
rect 92532 90352 92538 90364
rect 257430 90352 257436 90364
rect 92532 90324 257436 90352
rect 92532 90312 92538 90324
rect 257430 90312 257436 90324
rect 257488 90312 257494 90364
rect 336274 90312 336280 90364
rect 336332 90352 336338 90364
rect 556154 90352 556160 90364
rect 336332 90324 556160 90352
rect 336332 90312 336338 90324
rect 556154 90312 556160 90324
rect 556212 90312 556218 90364
rect 231854 89224 231860 89276
rect 231912 89264 231918 89276
rect 282086 89264 282092 89276
rect 231912 89236 282092 89264
rect 231912 89224 231918 89236
rect 282086 89224 282092 89236
rect 282144 89224 282150 89276
rect 301406 89224 301412 89276
rect 301464 89264 301470 89276
rect 347774 89264 347780 89276
rect 301464 89236 347780 89264
rect 301464 89224 301470 89236
rect 347774 89224 347780 89236
rect 347832 89224 347838 89276
rect 191834 89156 191840 89208
rect 191892 89196 191898 89208
rect 275554 89196 275560 89208
rect 191892 89168 275560 89196
rect 191892 89156 191898 89168
rect 275554 89156 275560 89168
rect 275612 89156 275618 89208
rect 305362 89156 305368 89208
rect 305420 89196 305426 89208
rect 371234 89196 371240 89208
rect 305420 89168 371240 89196
rect 305420 89156 305426 89168
rect 371234 89156 371240 89168
rect 371292 89156 371298 89208
rect 136634 89088 136640 89140
rect 136692 89128 136698 89140
rect 266354 89128 266360 89140
rect 136692 89100 266360 89128
rect 136692 89088 136698 89100
rect 266354 89088 266360 89100
rect 266412 89088 266418 89140
rect 315298 89088 315304 89140
rect 315356 89128 315362 89140
rect 411254 89128 411260 89140
rect 315356 89100 411260 89128
rect 315356 89088 315362 89100
rect 411254 89088 411260 89100
rect 411312 89088 411318 89140
rect 97994 89020 98000 89072
rect 98052 89060 98058 89072
rect 259914 89060 259920 89072
rect 98052 89032 259920 89060
rect 98052 89020 98058 89032
rect 259914 89020 259920 89032
rect 259972 89020 259978 89072
rect 339034 89020 339040 89072
rect 339092 89060 339098 89072
rect 494054 89060 494060 89072
rect 339092 89032 494060 89060
rect 339092 89020 339098 89032
rect 494054 89020 494060 89032
rect 494112 89020 494118 89072
rect 80054 88952 80060 89004
rect 80112 88992 80118 89004
rect 256786 88992 256792 89004
rect 80112 88964 256792 88992
rect 80112 88952 80118 88964
rect 256786 88952 256792 88964
rect 256844 88952 256850 89004
rect 329834 88952 329840 89004
rect 329892 88992 329898 89004
rect 517514 88992 517520 89004
rect 329892 88964 517520 88992
rect 329892 88952 329898 88964
rect 517514 88952 517520 88964
rect 517572 88952 517578 89004
rect 3326 88272 3332 88324
rect 3384 88312 3390 88324
rect 230106 88312 230112 88324
rect 3384 88284 230112 88312
rect 3384 88272 3390 88284
rect 230106 88272 230112 88284
rect 230164 88272 230170 88324
rect 354490 88272 354496 88324
rect 354548 88312 354554 88324
rect 580166 88312 580172 88324
rect 354548 88284 580172 88312
rect 354548 88272 354554 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 245838 87864 245844 87916
rect 245896 87904 245902 87916
rect 284386 87904 284392 87916
rect 245896 87876 284392 87904
rect 245896 87864 245902 87876
rect 284386 87864 284392 87876
rect 284444 87864 284450 87916
rect 223574 87796 223580 87848
rect 223632 87836 223638 87848
rect 280706 87836 280712 87848
rect 223632 87808 280712 87836
rect 223632 87796 223638 87808
rect 280706 87796 280712 87808
rect 280764 87796 280770 87848
rect 302050 87796 302056 87848
rect 302108 87836 302114 87848
rect 351914 87836 351920 87848
rect 302108 87808 351920 87836
rect 302108 87796 302114 87808
rect 351914 87796 351920 87808
rect 351972 87796 351978 87848
rect 208394 87728 208400 87780
rect 208452 87768 208458 87780
rect 278314 87768 278320 87780
rect 208452 87740 278320 87768
rect 208452 87728 208458 87740
rect 278314 87728 278320 87740
rect 278372 87728 278378 87780
rect 305914 87728 305920 87780
rect 305972 87768 305978 87780
rect 373994 87768 374000 87780
rect 305972 87740 374000 87768
rect 305972 87728 305978 87740
rect 373994 87728 374000 87740
rect 374052 87728 374058 87780
rect 187694 87660 187700 87712
rect 187752 87700 187758 87712
rect 272518 87700 272524 87712
rect 187752 87672 272524 87700
rect 187752 87660 187758 87672
rect 272518 87660 272524 87672
rect 272576 87660 272582 87712
rect 308306 87660 308312 87712
rect 308364 87700 308370 87712
rect 389174 87700 389180 87712
rect 308364 87672 389180 87700
rect 308364 87660 308370 87672
rect 389174 87660 389180 87672
rect 389232 87660 389238 87712
rect 115934 87592 115940 87644
rect 115992 87632 115998 87644
rect 262858 87632 262864 87644
rect 115992 87604 262864 87632
rect 115992 87592 115998 87604
rect 262858 87592 262864 87604
rect 262916 87592 262922 87644
rect 312538 87592 312544 87644
rect 312596 87632 312602 87644
rect 414014 87632 414020 87644
rect 312596 87604 414020 87632
rect 312596 87592 312602 87604
rect 414014 87592 414020 87604
rect 414072 87592 414078 87644
rect 235994 86436 236000 86488
rect 236052 86476 236058 86488
rect 282730 86476 282736 86488
rect 236052 86448 282736 86476
rect 236052 86436 236058 86448
rect 282730 86436 282736 86448
rect 282788 86436 282794 86488
rect 304810 86436 304816 86488
rect 304868 86476 304874 86488
rect 368474 86476 368480 86488
rect 304868 86448 368480 86476
rect 304868 86436 304874 86448
rect 368474 86436 368480 86448
rect 368532 86436 368538 86488
rect 197354 86368 197360 86420
rect 197412 86408 197418 86420
rect 276290 86408 276296 86420
rect 197412 86380 276296 86408
rect 197412 86368 197418 86380
rect 276290 86368 276296 86380
rect 276348 86368 276354 86420
rect 307754 86368 307760 86420
rect 307812 86408 307818 86420
rect 385034 86408 385040 86420
rect 307812 86380 385040 86408
rect 307812 86368 307818 86380
rect 385034 86368 385040 86380
rect 385092 86368 385098 86420
rect 139394 86300 139400 86352
rect 139452 86340 139458 86352
rect 264238 86340 264244 86352
rect 139452 86312 264244 86340
rect 139452 86300 139458 86312
rect 264238 86300 264244 86312
rect 264296 86300 264302 86352
rect 310882 86300 310888 86352
rect 310940 86340 310946 86352
rect 404354 86340 404360 86352
rect 310940 86312 404360 86340
rect 310940 86300 310946 86312
rect 404354 86300 404360 86312
rect 404412 86300 404418 86352
rect 89714 86232 89720 86284
rect 89772 86272 89778 86284
rect 255958 86272 255964 86284
rect 89772 86244 255964 86272
rect 89772 86232 89778 86244
rect 255958 86232 255964 86244
rect 256016 86232 256022 86284
rect 327994 86232 328000 86284
rect 328052 86272 328058 86284
rect 506474 86272 506480 86284
rect 328052 86244 506480 86272
rect 328052 86232 328058 86244
rect 506474 86232 506480 86244
rect 506532 86232 506538 86284
rect 230474 85076 230480 85128
rect 230532 85116 230538 85128
rect 281810 85116 281816 85128
rect 230532 85088 281816 85116
rect 230532 85076 230538 85088
rect 281810 85076 281816 85088
rect 281868 85076 281874 85128
rect 202874 85008 202880 85060
rect 202932 85048 202938 85060
rect 273990 85048 273996 85060
rect 202932 85020 273996 85048
rect 202932 85008 202938 85020
rect 273990 85008 273996 85020
rect 274048 85008 274054 85060
rect 306466 85008 306472 85060
rect 306524 85048 306530 85060
rect 378134 85048 378140 85060
rect 306524 85020 378140 85048
rect 306524 85008 306530 85020
rect 378134 85008 378140 85020
rect 378192 85008 378198 85060
rect 149054 84940 149060 84992
rect 149112 84980 149118 84992
rect 268378 84980 268384 84992
rect 149112 84952 268384 84980
rect 149112 84940 149118 84952
rect 268378 84940 268384 84952
rect 268436 84940 268442 84992
rect 312170 84940 312176 84992
rect 312228 84980 312234 84992
rect 412634 84980 412640 84992
rect 312228 84952 412640 84980
rect 312228 84940 312234 84952
rect 412634 84940 412640 84952
rect 412692 84940 412698 84992
rect 88334 84872 88340 84924
rect 88392 84912 88398 84924
rect 258258 84912 258264 84924
rect 88392 84884 258264 84912
rect 88392 84872 88398 84884
rect 258258 84872 258264 84884
rect 258316 84872 258322 84924
rect 314746 84872 314752 84924
rect 314804 84912 314810 84924
rect 427814 84912 427820 84924
rect 314804 84884 427820 84912
rect 314804 84872 314810 84884
rect 427814 84872 427820 84884
rect 427872 84872 427878 84924
rect 30374 84804 30380 84856
rect 30432 84844 30438 84856
rect 247678 84844 247684 84856
rect 30432 84816 247684 84844
rect 30432 84804 30438 84816
rect 247678 84804 247684 84816
rect 247736 84804 247742 84856
rect 328546 84804 328552 84856
rect 328604 84844 328610 84856
rect 510614 84844 510620 84856
rect 328604 84816 510620 84844
rect 328604 84804 328610 84816
rect 510614 84804 510620 84816
rect 510672 84804 510678 84856
rect 240134 83716 240140 83768
rect 240192 83756 240198 83768
rect 283190 83756 283196 83768
rect 240192 83728 283196 83756
rect 240192 83716 240198 83728
rect 283190 83716 283196 83728
rect 283248 83716 283254 83768
rect 215294 83648 215300 83700
rect 215352 83688 215358 83700
rect 279326 83688 279332 83700
rect 215352 83660 279332 83688
rect 215352 83648 215358 83660
rect 279326 83648 279332 83660
rect 279384 83648 279390 83700
rect 306926 83648 306932 83700
rect 306984 83688 306990 83700
rect 380894 83688 380900 83700
rect 306984 83660 380900 83688
rect 306984 83648 306990 83660
rect 380894 83648 380900 83660
rect 380952 83648 380958 83700
rect 158714 83580 158720 83632
rect 158772 83620 158778 83632
rect 269942 83620 269948 83632
rect 158772 83592 269948 83620
rect 158772 83580 158778 83592
rect 269942 83580 269948 83592
rect 270000 83580 270006 83632
rect 318058 83580 318064 83632
rect 318116 83620 318122 83632
rect 440326 83620 440332 83632
rect 318116 83592 440332 83620
rect 318116 83580 318122 83592
rect 440326 83580 440332 83592
rect 440384 83580 440390 83632
rect 70394 83512 70400 83564
rect 70452 83552 70458 83564
rect 255038 83552 255044 83564
rect 70452 83524 255044 83552
rect 70452 83512 70458 83524
rect 255038 83512 255044 83524
rect 255096 83512 255102 83564
rect 320358 83512 320364 83564
rect 320416 83552 320422 83564
rect 462406 83552 462412 83564
rect 320416 83524 462412 83552
rect 320416 83512 320422 83524
rect 462406 83512 462412 83524
rect 462464 83512 462470 83564
rect 53834 83444 53840 83496
rect 53892 83484 53898 83496
rect 252554 83484 252560 83496
rect 53892 83456 252560 83484
rect 53892 83444 53898 83456
rect 252554 83444 252560 83456
rect 252612 83444 252618 83496
rect 294414 83444 294420 83496
rect 294472 83484 294478 83496
rect 306374 83484 306380 83496
rect 294472 83456 306380 83484
rect 294472 83444 294478 83456
rect 306374 83444 306380 83456
rect 306432 83444 306438 83496
rect 329006 83444 329012 83496
rect 329064 83484 329070 83496
rect 513374 83484 513380 83496
rect 329064 83456 513380 83484
rect 329064 83444 329070 83456
rect 513374 83444 513380 83456
rect 513432 83444 513438 83496
rect 222194 82288 222200 82340
rect 222252 82328 222258 82340
rect 279602 82328 279608 82340
rect 222252 82300 279608 82328
rect 222252 82288 222258 82300
rect 279602 82288 279608 82300
rect 279660 82288 279666 82340
rect 301774 82288 301780 82340
rect 301832 82328 301838 82340
rect 350534 82328 350540 82340
rect 301832 82300 350540 82328
rect 301832 82288 301838 82300
rect 350534 82288 350540 82300
rect 350592 82288 350598 82340
rect 165614 82220 165620 82272
rect 165672 82260 165678 82272
rect 271046 82260 271052 82272
rect 165672 82232 271052 82260
rect 165672 82220 165678 82232
rect 271046 82220 271052 82232
rect 271104 82220 271110 82272
rect 309134 82220 309140 82272
rect 309192 82260 309198 82272
rect 394694 82260 394700 82272
rect 309192 82232 394700 82260
rect 309192 82220 309198 82232
rect 394694 82220 394700 82232
rect 394752 82220 394758 82272
rect 138014 82152 138020 82204
rect 138072 82192 138078 82204
rect 266446 82192 266452 82204
rect 138072 82164 266452 82192
rect 138072 82152 138078 82164
rect 266446 82152 266452 82164
rect 266504 82152 266510 82204
rect 329558 82152 329564 82204
rect 329616 82192 329622 82204
rect 517606 82192 517612 82204
rect 329616 82164 517612 82192
rect 329616 82152 329622 82164
rect 517606 82152 517612 82164
rect 517664 82152 517670 82204
rect 42794 82084 42800 82136
rect 42852 82124 42858 82136
rect 250622 82124 250628 82136
rect 42852 82096 250628 82124
rect 42852 82084 42858 82096
rect 250622 82084 250628 82096
rect 250680 82084 250686 82136
rect 323946 82084 323952 82136
rect 324004 82124 324010 82136
rect 328454 82124 328460 82136
rect 324004 82096 328460 82124
rect 324004 82084 324010 82096
rect 328454 82084 328460 82096
rect 328512 82084 328518 82136
rect 333054 82084 333060 82136
rect 333112 82124 333118 82136
rect 538214 82124 538220 82136
rect 333112 82096 538220 82124
rect 333112 82084 333118 82096
rect 538214 82084 538220 82096
rect 538272 82084 538278 82136
rect 220814 80860 220820 80912
rect 220872 80900 220878 80912
rect 280338 80900 280344 80912
rect 220872 80872 280344 80900
rect 220872 80860 220878 80872
rect 280338 80860 280344 80872
rect 280396 80860 280402 80912
rect 300118 80860 300124 80912
rect 300176 80900 300182 80912
rect 340966 80900 340972 80912
rect 300176 80872 340972 80900
rect 300176 80860 300182 80872
rect 340966 80860 340972 80872
rect 341024 80860 341030 80912
rect 190454 80792 190460 80844
rect 190512 80832 190518 80844
rect 275186 80832 275192 80844
rect 190512 80804 275192 80832
rect 190512 80792 190518 80804
rect 275186 80792 275192 80804
rect 275244 80792 275250 80844
rect 307478 80792 307484 80844
rect 307536 80832 307542 80844
rect 385126 80832 385132 80844
rect 307536 80804 385132 80832
rect 307536 80792 307542 80804
rect 385126 80792 385132 80804
rect 385184 80792 385190 80844
rect 142154 80724 142160 80776
rect 142212 80764 142218 80776
rect 265618 80764 265624 80776
rect 142212 80736 265624 80764
rect 142212 80724 142218 80736
rect 265618 80724 265624 80736
rect 265676 80724 265682 80776
rect 338942 80724 338948 80776
rect 339000 80764 339006 80776
rect 520274 80764 520280 80776
rect 339000 80736 520280 80764
rect 339000 80724 339006 80736
rect 520274 80724 520280 80736
rect 520332 80724 520338 80776
rect 120074 80656 120080 80708
rect 120132 80696 120138 80708
rect 263318 80696 263324 80708
rect 120132 80668 263324 80696
rect 120132 80656 120138 80668
rect 263318 80656 263324 80668
rect 263376 80656 263382 80708
rect 330294 80656 330300 80708
rect 330352 80696 330358 80708
rect 521654 80696 521660 80708
rect 330352 80668 521660 80696
rect 330352 80656 330358 80668
rect 521654 80656 521660 80668
rect 521712 80656 521718 80708
rect 302234 79500 302240 79552
rect 302292 79540 302298 79552
rect 352006 79540 352012 79552
rect 302292 79512 352012 79540
rect 302292 79500 302298 79512
rect 352006 79500 352012 79512
rect 352064 79500 352070 79552
rect 202966 79432 202972 79484
rect 203024 79472 203030 79484
rect 277670 79472 277676 79484
rect 203024 79444 277676 79472
rect 203024 79432 203030 79444
rect 277670 79432 277676 79444
rect 277728 79432 277734 79484
rect 311342 79432 311348 79484
rect 311400 79472 311406 79484
rect 407114 79472 407120 79484
rect 311400 79444 407120 79472
rect 311400 79432 311406 79444
rect 407114 79432 407120 79444
rect 407172 79432 407178 79484
rect 146294 79364 146300 79416
rect 146352 79404 146358 79416
rect 267734 79404 267740 79416
rect 146352 79376 267740 79404
rect 146352 79364 146358 79376
rect 267734 79364 267740 79376
rect 267792 79364 267798 79416
rect 313274 79364 313280 79416
rect 313332 79404 313338 79416
rect 418154 79404 418160 79416
rect 313332 79376 418160 79404
rect 313332 79364 313338 79376
rect 418154 79364 418160 79376
rect 418212 79364 418218 79416
rect 96614 79296 96620 79348
rect 96672 79336 96678 79348
rect 259454 79336 259460 79348
rect 96672 79308 259460 79336
rect 96672 79296 96678 79308
rect 259454 79296 259460 79308
rect 259512 79296 259518 79348
rect 331766 79296 331772 79348
rect 331824 79336 331830 79348
rect 529934 79336 529940 79348
rect 331824 79308 529940 79336
rect 331824 79296 331830 79308
rect 529934 79296 529940 79308
rect 529992 79296 529998 79348
rect 207014 78140 207020 78192
rect 207072 78180 207078 78192
rect 277946 78180 277952 78192
rect 207072 78152 277952 78180
rect 207072 78140 207078 78152
rect 277946 78140 277952 78152
rect 278004 78140 278010 78192
rect 303246 78140 303252 78192
rect 303304 78180 303310 78192
rect 358814 78180 358820 78192
rect 303304 78152 358820 78180
rect 303304 78140 303310 78152
rect 358814 78140 358820 78152
rect 358872 78140 358878 78192
rect 153194 78072 153200 78124
rect 153252 78112 153258 78124
rect 268838 78112 268844 78124
rect 153252 78084 268844 78112
rect 153252 78072 153258 78084
rect 268838 78072 268844 78084
rect 268896 78072 268902 78124
rect 312998 78072 313004 78124
rect 313056 78112 313062 78124
rect 418246 78112 418252 78124
rect 313056 78084 418252 78112
rect 313056 78072 313062 78084
rect 418246 78072 418252 78084
rect 418304 78072 418310 78124
rect 99374 78004 99380 78056
rect 99432 78044 99438 78056
rect 260006 78044 260012 78056
rect 99432 78016 260012 78044
rect 99432 78004 99438 78016
rect 260006 78004 260012 78016
rect 260064 78004 260070 78056
rect 317046 78004 317052 78056
rect 317104 78044 317110 78056
rect 441614 78044 441620 78056
rect 317104 78016 441620 78044
rect 317104 78004 317110 78016
rect 441614 78004 441620 78016
rect 441672 78004 441678 78056
rect 78674 77936 78680 77988
rect 78732 77976 78738 77988
rect 256510 77976 256516 77988
rect 78732 77948 256516 77976
rect 78732 77936 78738 77948
rect 256510 77936 256516 77948
rect 256568 77936 256574 77988
rect 332318 77936 332324 77988
rect 332376 77976 332382 77988
rect 534074 77976 534080 77988
rect 332376 77948 534080 77976
rect 332376 77936 332382 77948
rect 534074 77936 534080 77948
rect 534132 77936 534138 77988
rect 226334 76712 226340 76764
rect 226392 76752 226398 76764
rect 281166 76752 281172 76764
rect 226392 76724 281172 76752
rect 226392 76712 226398 76724
rect 281166 76712 281172 76724
rect 281224 76712 281230 76764
rect 300486 76712 300492 76764
rect 300544 76752 300550 76764
rect 342254 76752 342260 76764
rect 300544 76724 342260 76752
rect 300544 76712 300550 76724
rect 342254 76712 342260 76724
rect 342312 76712 342318 76764
rect 162854 76644 162860 76696
rect 162912 76684 162918 76696
rect 270494 76684 270500 76696
rect 162912 76656 270500 76684
rect 162912 76644 162918 76656
rect 270494 76644 270500 76656
rect 270552 76644 270558 76696
rect 305454 76644 305460 76696
rect 305512 76684 305518 76696
rect 372614 76684 372620 76696
rect 305512 76656 372620 76684
rect 305512 76644 305518 76656
rect 372614 76644 372620 76656
rect 372672 76644 372678 76696
rect 82814 76576 82820 76628
rect 82872 76616 82878 76628
rect 257246 76616 257252 76628
rect 82872 76588 257252 76616
rect 82872 76576 82878 76588
rect 257246 76576 257252 76588
rect 257304 76576 257310 76628
rect 326338 76576 326344 76628
rect 326396 76616 326402 76628
rect 437474 76616 437480 76628
rect 326396 76588 437480 76616
rect 326396 76576 326402 76588
rect 437474 76576 437480 76588
rect 437532 76576 437538 76628
rect 35894 76508 35900 76560
rect 35952 76548 35958 76560
rect 249334 76548 249340 76560
rect 35952 76520 249340 76548
rect 35952 76508 35958 76520
rect 249334 76508 249340 76520
rect 249392 76508 249398 76560
rect 337470 76508 337476 76560
rect 337528 76548 337534 76560
rect 546494 76548 546500 76560
rect 337528 76520 546500 76548
rect 337528 76508 337534 76520
rect 546494 76508 546500 76520
rect 546552 76508 546558 76560
rect 354398 75828 354404 75880
rect 354456 75868 354462 75880
rect 580166 75868 580172 75880
rect 354456 75840 580172 75868
rect 354456 75828 354462 75840
rect 580166 75828 580172 75840
rect 580224 75828 580230 75880
rect 236086 75352 236092 75404
rect 236144 75392 236150 75404
rect 283006 75392 283012 75404
rect 236144 75364 283012 75392
rect 236144 75352 236150 75364
rect 283006 75352 283012 75364
rect 283064 75352 283070 75404
rect 169846 75284 169852 75336
rect 169904 75324 169910 75336
rect 271138 75324 271144 75336
rect 169904 75296 271144 75324
rect 169904 75284 169910 75296
rect 271138 75284 271144 75296
rect 271196 75284 271202 75336
rect 301590 75284 301596 75336
rect 301648 75324 301654 75336
rect 349154 75324 349160 75336
rect 301648 75296 349160 75324
rect 301648 75284 301654 75296
rect 349154 75284 349160 75296
rect 349212 75284 349218 75336
rect 103514 75216 103520 75268
rect 103572 75256 103578 75268
rect 261018 75256 261024 75268
rect 103572 75228 261024 75256
rect 103572 75216 103578 75228
rect 261018 75216 261024 75228
rect 261076 75216 261082 75268
rect 310974 75216 310980 75268
rect 311032 75256 311038 75268
rect 405734 75256 405740 75268
rect 311032 75228 405740 75256
rect 311032 75216 311038 75228
rect 405734 75216 405740 75228
rect 405792 75216 405798 75268
rect 26234 75148 26240 75200
rect 26292 75188 26298 75200
rect 246390 75188 246396 75200
rect 26292 75160 246396 75188
rect 26292 75148 26298 75160
rect 246390 75148 246396 75160
rect 246448 75148 246454 75200
rect 314102 75148 314108 75200
rect 314160 75188 314166 75200
rect 423674 75188 423680 75200
rect 314160 75160 423680 75188
rect 314160 75148 314166 75160
rect 423674 75148 423680 75160
rect 423732 75148 423738 75200
rect 3326 74468 3332 74520
rect 3384 74508 3390 74520
rect 230014 74508 230020 74520
rect 3384 74480 230020 74508
rect 3384 74468 3390 74480
rect 230014 74468 230020 74480
rect 230072 74468 230078 74520
rect 225046 73924 225052 73976
rect 225104 73964 225110 73976
rect 280798 73964 280804 73976
rect 225104 73936 280804 73964
rect 225104 73924 225110 73936
rect 280798 73924 280804 73936
rect 280856 73924 280862 73976
rect 304994 73924 305000 73976
rect 305052 73964 305058 73976
rect 368566 73964 368572 73976
rect 305052 73936 368572 73964
rect 305052 73924 305058 73936
rect 368566 73924 368572 73936
rect 368624 73924 368630 73976
rect 200114 73856 200120 73908
rect 200172 73896 200178 73908
rect 276842 73896 276848 73908
rect 200172 73868 276848 73896
rect 200172 73856 200178 73868
rect 276842 73856 276848 73868
rect 276900 73856 276906 73908
rect 321554 73856 321560 73908
rect 321612 73896 321618 73908
rect 467926 73896 467932 73908
rect 321612 73868 467932 73896
rect 321612 73856 321618 73868
rect 467926 73856 467932 73868
rect 467984 73856 467990 73908
rect 91094 73788 91100 73840
rect 91152 73828 91158 73840
rect 258626 73828 258632 73840
rect 91152 73800 258632 73828
rect 91152 73788 91158 73800
rect 258626 73788 258632 73800
rect 258684 73788 258690 73840
rect 276014 73788 276020 73840
rect 276072 73828 276078 73840
rect 289446 73828 289452 73840
rect 276072 73800 289452 73828
rect 276072 73788 276078 73800
rect 289446 73788 289452 73800
rect 289504 73788 289510 73840
rect 335078 73788 335084 73840
rect 335136 73828 335142 73840
rect 549898 73828 549904 73840
rect 335136 73800 549904 73828
rect 335136 73788 335142 73800
rect 549898 73788 549904 73800
rect 549956 73788 549962 73840
rect 302694 72632 302700 72684
rect 302752 72672 302758 72684
rect 356054 72672 356060 72684
rect 302752 72644 356060 72672
rect 302752 72632 302758 72644
rect 356054 72632 356060 72644
rect 356112 72632 356118 72684
rect 176654 72564 176660 72616
rect 176712 72604 176718 72616
rect 272886 72604 272892 72616
rect 176712 72576 272892 72604
rect 176712 72564 176718 72576
rect 272886 72564 272892 72576
rect 272944 72564 272950 72616
rect 308766 72564 308772 72616
rect 308824 72604 308830 72616
rect 391934 72604 391940 72616
rect 308824 72576 391940 72604
rect 308824 72564 308830 72576
rect 391934 72564 391940 72576
rect 391992 72564 391998 72616
rect 153286 72496 153292 72548
rect 153344 72536 153350 72548
rect 269298 72536 269304 72548
rect 153344 72508 269304 72536
rect 153344 72496 153350 72508
rect 269298 72496 269304 72508
rect 269356 72496 269362 72548
rect 324406 72496 324412 72548
rect 324464 72536 324470 72548
rect 485774 72536 485780 72548
rect 324464 72508 485780 72536
rect 324464 72496 324470 72508
rect 485774 72496 485780 72508
rect 485832 72496 485838 72548
rect 46934 72428 46940 72480
rect 46992 72468 46998 72480
rect 251174 72468 251180 72480
rect 46992 72440 251180 72468
rect 46992 72428 46998 72440
rect 251174 72428 251180 72440
rect 251232 72428 251238 72480
rect 298830 72428 298836 72480
rect 298888 72468 298894 72480
rect 332594 72468 332600 72480
rect 298888 72440 332600 72468
rect 298888 72428 298894 72440
rect 332594 72428 332600 72440
rect 332652 72428 332658 72480
rect 337378 72428 337384 72480
rect 337436 72468 337442 72480
rect 553394 72468 553400 72480
rect 337436 72440 553400 72468
rect 337436 72428 337442 72440
rect 553394 72428 553400 72440
rect 553452 72428 553458 72480
rect 197446 71136 197452 71188
rect 197504 71176 197510 71188
rect 276382 71176 276388 71188
rect 197504 71148 276388 71176
rect 197504 71136 197510 71148
rect 276382 71136 276388 71148
rect 276440 71136 276446 71188
rect 309686 71136 309692 71188
rect 309744 71176 309750 71188
rect 397454 71176 397460 71188
rect 309744 71148 397460 71176
rect 309744 71136 309750 71148
rect 397454 71136 397460 71148
rect 397512 71136 397518 71188
rect 180794 71068 180800 71120
rect 180852 71108 180858 71120
rect 273530 71108 273536 71120
rect 180852 71080 273536 71108
rect 180852 71068 180858 71080
rect 273530 71068 273536 71080
rect 273588 71068 273594 71120
rect 316494 71068 316500 71120
rect 316552 71108 316558 71120
rect 438854 71108 438860 71120
rect 316552 71080 438860 71108
rect 316552 71068 316558 71080
rect 438854 71068 438860 71080
rect 438912 71068 438918 71120
rect 109034 71000 109040 71052
rect 109092 71040 109098 71052
rect 261662 71040 261668 71052
rect 109092 71012 261668 71040
rect 109092 71000 109098 71012
rect 261662 71000 261668 71012
rect 261720 71000 261726 71052
rect 273254 71000 273260 71052
rect 273312 71040 273318 71052
rect 288986 71040 288992 71052
rect 273312 71012 288992 71040
rect 273312 71000 273318 71012
rect 288986 71000 288992 71012
rect 289044 71000 289050 71052
rect 319622 71000 319628 71052
rect 319680 71040 319686 71052
rect 456886 71040 456892 71052
rect 319680 71012 456892 71040
rect 319680 71000 319686 71012
rect 456886 71000 456892 71012
rect 456944 71000 456950 71052
rect 201494 69776 201500 69828
rect 201552 69816 201558 69828
rect 276934 69816 276940 69828
rect 201552 69788 276940 69816
rect 201552 69776 201558 69788
rect 276934 69776 276940 69788
rect 276992 69776 276998 69828
rect 310238 69776 310244 69828
rect 310296 69816 310302 69828
rect 401594 69816 401600 69828
rect 310296 69788 401600 69816
rect 310296 69776 310302 69788
rect 401594 69776 401600 69788
rect 401652 69776 401658 69828
rect 183554 69708 183560 69760
rect 183612 69748 183618 69760
rect 273622 69748 273628 69760
rect 183612 69720 273628 69748
rect 183612 69708 183618 69720
rect 273622 69708 273628 69720
rect 273680 69708 273686 69760
rect 320174 69708 320180 69760
rect 320232 69748 320238 69760
rect 460934 69748 460940 69760
rect 320232 69720 460940 69748
rect 320232 69708 320238 69720
rect 460934 69708 460940 69720
rect 460992 69708 460998 69760
rect 113174 69640 113180 69692
rect 113232 69680 113238 69692
rect 260098 69680 260104 69692
rect 113232 69652 260104 69680
rect 113232 69640 113238 69652
rect 260098 69640 260104 69652
rect 260156 69640 260162 69692
rect 294966 69640 294972 69692
rect 295024 69680 295030 69692
rect 309134 69680 309140 69692
rect 295024 69652 309140 69680
rect 295024 69640 295030 69652
rect 309134 69640 309140 69652
rect 309192 69640 309198 69692
rect 322750 69640 322756 69692
rect 322808 69680 322814 69692
rect 476114 69680 476120 69692
rect 322808 69652 476120 69680
rect 322808 69640 322814 69652
rect 476114 69640 476120 69652
rect 476172 69640 476178 69692
rect 234614 68484 234620 68536
rect 234672 68524 234678 68536
rect 282454 68524 282460 68536
rect 234672 68496 282460 68524
rect 234672 68484 234678 68496
rect 282454 68484 282460 68496
rect 282512 68484 282518 68536
rect 186314 68416 186320 68468
rect 186372 68456 186378 68468
rect 274910 68456 274916 68468
rect 186372 68428 274916 68456
rect 186372 68416 186378 68428
rect 274910 68416 274916 68428
rect 274968 68416 274974 68468
rect 315206 68416 315212 68468
rect 315264 68456 315270 68468
rect 430574 68456 430580 68468
rect 315264 68428 430580 68456
rect 315264 68416 315270 68428
rect 430574 68416 430580 68428
rect 430632 68416 430638 68468
rect 86954 68348 86960 68400
rect 87012 68388 87018 68400
rect 257798 68388 257804 68400
rect 87012 68360 257804 68388
rect 87012 68348 87018 68360
rect 257798 68348 257804 68360
rect 257856 68348 257862 68400
rect 324774 68348 324780 68400
rect 324832 68388 324838 68400
rect 488534 68388 488540 68400
rect 324832 68360 488540 68388
rect 324832 68348 324838 68360
rect 488534 68348 488540 68360
rect 488592 68348 488598 68400
rect 57974 68280 57980 68332
rect 58032 68320 58038 68332
rect 253014 68320 253020 68332
rect 58032 68292 253020 68320
rect 58032 68280 58038 68292
rect 253014 68280 253020 68292
rect 253072 68280 253078 68332
rect 332778 68280 332784 68332
rect 332836 68320 332842 68332
rect 535454 68320 535460 68332
rect 332836 68292 535460 68320
rect 332836 68280 332842 68292
rect 535454 68280 535460 68292
rect 535512 68280 535518 68332
rect 193214 66988 193220 67040
rect 193272 67028 193278 67040
rect 275646 67028 275652 67040
rect 193272 67000 275652 67028
rect 193272 66988 193278 67000
rect 275646 66988 275652 67000
rect 275704 66988 275710 67040
rect 303982 66988 303988 67040
rect 304040 67028 304046 67040
rect 363046 67028 363052 67040
rect 304040 67000 363052 67028
rect 304040 66988 304046 67000
rect 363046 66988 363052 67000
rect 363104 66988 363110 67040
rect 114554 66920 114560 66972
rect 114612 66960 114618 66972
rect 262490 66960 262496 66972
rect 114612 66932 262496 66960
rect 114612 66920 114618 66932
rect 262490 66920 262496 66932
rect 262548 66920 262554 66972
rect 315758 66920 315764 66972
rect 315816 66960 315822 66972
rect 434806 66960 434812 66972
rect 315816 66932 434812 66960
rect 315816 66920 315822 66932
rect 434806 66920 434812 66932
rect 434864 66920 434870 66972
rect 20714 66852 20720 66904
rect 20772 66892 20778 66904
rect 243630 66892 243636 66904
rect 20772 66864 243636 66892
rect 20772 66852 20778 66864
rect 243630 66852 243636 66864
rect 243688 66852 243694 66904
rect 325878 66852 325884 66904
rect 325936 66892 325942 66904
rect 495434 66892 495440 66904
rect 325936 66864 495440 66892
rect 325936 66852 325942 66864
rect 495434 66852 495440 66864
rect 495492 66852 495498 66904
rect 214006 65628 214012 65680
rect 214064 65668 214070 65680
rect 279142 65668 279148 65680
rect 214064 65640 279148 65668
rect 214064 65628 214070 65640
rect 279142 65628 279148 65640
rect 279200 65628 279206 65680
rect 309502 65628 309508 65680
rect 309560 65668 309566 65680
rect 396074 65668 396080 65680
rect 309560 65640 396080 65668
rect 309560 65628 309566 65640
rect 396074 65628 396080 65640
rect 396132 65628 396138 65680
rect 140774 65560 140780 65612
rect 140832 65600 140838 65612
rect 266814 65600 266820 65612
rect 140832 65572 266820 65600
rect 140832 65560 140838 65572
rect 266814 65560 266820 65572
rect 266872 65560 266878 65612
rect 317414 65560 317420 65612
rect 317472 65600 317478 65612
rect 444374 65600 444380 65612
rect 317472 65572 444380 65600
rect 317472 65560 317478 65572
rect 444374 65560 444380 65572
rect 444432 65560 444438 65612
rect 59354 65492 59360 65544
rect 59412 65532 59418 65544
rect 253382 65532 253388 65544
rect 59412 65504 253388 65532
rect 59412 65492 59418 65504
rect 253382 65492 253388 65504
rect 253440 65492 253446 65544
rect 327534 65492 327540 65544
rect 327592 65532 327598 65544
rect 505094 65532 505100 65544
rect 327592 65504 505100 65532
rect 327592 65492 327598 65504
rect 505094 65492 505100 65504
rect 505152 65492 505158 65544
rect 209774 64268 209780 64320
rect 209832 64308 209838 64320
rect 278406 64308 278412 64320
rect 209832 64280 278412 64308
rect 209832 64268 209838 64280
rect 278406 64268 278412 64280
rect 278464 64268 278470 64320
rect 314470 64268 314476 64320
rect 314528 64308 314534 64320
rect 426434 64308 426440 64320
rect 314528 64280 426440 64308
rect 314528 64268 314534 64280
rect 426434 64268 426440 64280
rect 426492 64268 426498 64320
rect 161474 64200 161480 64252
rect 161532 64240 161538 64252
rect 270310 64240 270316 64252
rect 161532 64212 270316 64240
rect 161532 64200 161538 64212
rect 270310 64200 270316 64212
rect 270368 64200 270374 64252
rect 317966 64200 317972 64252
rect 318024 64240 318030 64252
rect 447134 64240 447140 64252
rect 318024 64212 447140 64240
rect 318024 64200 318030 64212
rect 447134 64200 447140 64212
rect 447192 64200 447198 64252
rect 49694 64132 49700 64184
rect 49752 64172 49758 64184
rect 251726 64172 251732 64184
rect 49752 64144 251732 64172
rect 49752 64132 49758 64144
rect 251726 64132 251732 64144
rect 251784 64132 251790 64184
rect 296806 64132 296812 64184
rect 296864 64172 296870 64184
rect 320174 64172 320180 64184
rect 296864 64144 320180 64172
rect 296864 64132 296870 64144
rect 320174 64132 320180 64144
rect 320232 64132 320238 64184
rect 330846 64132 330852 64184
rect 330904 64172 330910 64184
rect 524414 64172 524420 64184
rect 330904 64144 524420 64172
rect 330904 64132 330910 64144
rect 524414 64132 524420 64144
rect 524472 64132 524478 64184
rect 266446 62976 266452 63028
rect 266504 63016 266510 63028
rect 287790 63016 287796 63028
rect 266504 62988 287796 63016
rect 266504 62976 266510 62988
rect 287790 62976 287796 62988
rect 287848 62976 287854 63028
rect 312262 62908 312268 62960
rect 312320 62948 312326 62960
rect 412726 62948 412732 62960
rect 312320 62920 412732 62948
rect 312320 62908 312326 62920
rect 412726 62908 412732 62920
rect 412784 62908 412790 62960
rect 143534 62840 143540 62892
rect 143592 62880 143598 62892
rect 267366 62880 267372 62892
rect 143592 62852 267372 62880
rect 143592 62840 143598 62852
rect 267366 62840 267372 62852
rect 267424 62840 267430 62892
rect 318518 62840 318524 62892
rect 318576 62880 318582 62892
rect 451274 62880 451280 62892
rect 318576 62852 451280 62880
rect 318576 62840 318582 62852
rect 451274 62840 451280 62852
rect 451332 62840 451338 62892
rect 103606 62772 103612 62824
rect 103664 62812 103670 62824
rect 260558 62812 260564 62824
rect 103664 62784 260564 62812
rect 103664 62772 103670 62784
rect 260558 62772 260564 62784
rect 260616 62772 260622 62824
rect 296254 62772 296260 62824
rect 296312 62812 296318 62824
rect 317414 62812 317420 62824
rect 296312 62784 317420 62812
rect 296312 62772 296318 62784
rect 317414 62772 317420 62784
rect 317472 62772 317478 62824
rect 332686 62772 332692 62824
rect 332744 62812 332750 62824
rect 534166 62812 534172 62824
rect 332744 62784 534172 62812
rect 332744 62772 332750 62784
rect 534166 62772 534172 62784
rect 534224 62772 534230 62824
rect 354306 62024 354312 62076
rect 354364 62064 354370 62076
rect 580166 62064 580172 62076
rect 354364 62036 580172 62064
rect 354364 62024 354370 62036
rect 580166 62024 580172 62036
rect 580224 62024 580230 62076
rect 242894 61548 242900 61600
rect 242952 61588 242958 61600
rect 283926 61588 283932 61600
rect 242952 61560 283932 61588
rect 242952 61548 242958 61560
rect 283926 61548 283932 61560
rect 283984 61548 283990 61600
rect 171134 61480 171140 61532
rect 171192 61520 171198 61532
rect 272058 61520 272064 61532
rect 171192 61492 272064 61520
rect 171192 61480 171198 61492
rect 272058 61480 272064 61492
rect 272116 61480 272122 61532
rect 299474 61480 299480 61532
rect 299532 61520 299538 61532
rect 335354 61520 335360 61532
rect 299532 61492 335360 61520
rect 299532 61480 299538 61492
rect 335354 61480 335360 61492
rect 335412 61480 335418 61532
rect 122834 61412 122840 61464
rect 122892 61452 122898 61464
rect 263870 61452 263876 61464
rect 122892 61424 263876 61452
rect 122892 61412 122898 61424
rect 263870 61412 263876 61424
rect 263928 61412 263934 61464
rect 304350 61412 304356 61464
rect 304408 61452 304414 61464
rect 365714 61452 365720 61464
rect 304408 61424 365720 61452
rect 304408 61412 304414 61424
rect 365714 61412 365720 61424
rect 365772 61412 365778 61464
rect 35158 61344 35164 61396
rect 35216 61384 35222 61396
rect 248874 61384 248880 61396
rect 35216 61356 248880 61384
rect 35216 61344 35222 61356
rect 248874 61344 248880 61356
rect 248932 61344 248938 61396
rect 319254 61344 319260 61396
rect 319312 61384 319318 61396
rect 455414 61384 455420 61396
rect 319312 61356 455420 61384
rect 319312 61344 319318 61356
rect 455414 61344 455420 61356
rect 455472 61344 455478 61396
rect 313366 60120 313372 60172
rect 313424 60160 313430 60172
rect 419534 60160 419540 60172
rect 313424 60132 419540 60160
rect 313424 60120 313430 60132
rect 419534 60120 419540 60132
rect 419592 60120 419598 60172
rect 147674 60052 147680 60104
rect 147732 60092 147738 60104
rect 268010 60092 268016 60104
rect 147732 60064 268016 60092
rect 147732 60052 147738 60064
rect 268010 60052 268016 60064
rect 268068 60052 268074 60104
rect 320726 60052 320732 60104
rect 320784 60092 320790 60104
rect 463694 60092 463700 60104
rect 320784 60064 463700 60092
rect 320784 60052 320790 60064
rect 463694 60052 463700 60064
rect 463752 60052 463758 60104
rect 125594 59984 125600 60036
rect 125652 60024 125658 60036
rect 264422 60024 264428 60036
rect 125652 59996 264428 60024
rect 125652 59984 125658 59996
rect 264422 59984 264428 59996
rect 264480 59984 264486 60036
rect 295702 59984 295708 60036
rect 295760 60024 295766 60036
rect 313274 60024 313280 60036
rect 295760 59996 313280 60024
rect 295760 59984 295766 59996
rect 313274 59984 313280 59996
rect 313332 59984 313338 60036
rect 335814 59984 335820 60036
rect 335872 60024 335878 60036
rect 552658 60024 552664 60036
rect 335872 59996 552664 60024
rect 335872 59984 335878 59996
rect 552658 59984 552664 59996
rect 552716 59984 552722 60036
rect 306558 58760 306564 58812
rect 306616 58800 306622 58812
rect 379514 58800 379520 58812
rect 306616 58772 379520 58800
rect 306616 58760 306622 58772
rect 379514 58760 379520 58772
rect 379572 58760 379578 58812
rect 150434 58692 150440 58744
rect 150492 58732 150498 58744
rect 268470 58732 268476 58744
rect 150492 58704 268476 58732
rect 150492 58692 150498 58704
rect 268470 58692 268476 58704
rect 268528 58692 268534 58744
rect 322014 58692 322020 58744
rect 322072 58732 322078 58744
rect 471974 58732 471980 58744
rect 322072 58704 471980 58732
rect 322072 58692 322078 58704
rect 471974 58692 471980 58704
rect 472032 58692 472038 58744
rect 129734 58624 129740 58676
rect 129792 58664 129798 58676
rect 265066 58664 265072 58676
rect 129792 58636 265072 58664
rect 129792 58624 129798 58636
rect 265066 58624 265072 58636
rect 265124 58624 265130 58676
rect 327166 58624 327172 58676
rect 327224 58664 327230 58676
rect 502334 58664 502340 58676
rect 327224 58636 502340 58664
rect 327224 58624 327230 58636
rect 502334 58624 502340 58636
rect 502392 58624 502398 58676
rect 307110 57332 307116 57384
rect 307168 57372 307174 57384
rect 382274 57372 382280 57384
rect 307168 57344 382280 57372
rect 307168 57332 307174 57344
rect 382274 57332 382280 57344
rect 382332 57332 382338 57384
rect 157334 57264 157340 57316
rect 157392 57304 157398 57316
rect 269574 57304 269580 57316
rect 157392 57276 269580 57304
rect 157392 57264 157398 57276
rect 269574 57264 269580 57276
rect 269632 57264 269638 57316
rect 322566 57264 322572 57316
rect 322624 57304 322630 57316
rect 474734 57304 474740 57316
rect 322624 57276 474740 57304
rect 322624 57264 322630 57276
rect 474734 57264 474740 57276
rect 474792 57264 474798 57316
rect 132494 57196 132500 57248
rect 132552 57236 132558 57248
rect 265158 57236 265164 57248
rect 132552 57208 265164 57236
rect 132552 57196 132558 57208
rect 265158 57196 265164 57208
rect 265216 57196 265222 57248
rect 331030 57196 331036 57248
rect 331088 57236 331094 57248
rect 525794 57236 525800 57248
rect 331088 57208 525800 57236
rect 331088 57196 331094 57208
rect 525794 57196 525800 57208
rect 525852 57196 525858 57248
rect 309318 55972 309324 56024
rect 309376 56012 309382 56024
rect 396166 56012 396172 56024
rect 309376 55984 396172 56012
rect 309376 55972 309382 55984
rect 396166 55972 396172 55984
rect 396224 55972 396230 56024
rect 160094 55904 160100 55956
rect 160152 55944 160158 55956
rect 270126 55944 270132 55956
rect 160152 55916 270132 55944
rect 160152 55904 160158 55916
rect 270126 55904 270132 55916
rect 270184 55904 270190 55956
rect 323118 55904 323124 55956
rect 323176 55944 323182 55956
rect 478874 55944 478880 55956
rect 323176 55916 478880 55944
rect 323176 55904 323182 55916
rect 478874 55904 478880 55916
rect 478932 55904 478938 55956
rect 53926 55836 53932 55888
rect 53984 55876 53990 55888
rect 252278 55876 252284 55888
rect 53984 55848 252284 55876
rect 53984 55836 53990 55848
rect 252278 55836 252284 55848
rect 252336 55836 252342 55888
rect 334342 55836 334348 55888
rect 334400 55876 334406 55888
rect 545114 55876 545120 55888
rect 334400 55848 545120 55876
rect 334400 55836 334406 55848
rect 545114 55836 545120 55848
rect 545172 55836 545178 55888
rect 164234 54544 164240 54596
rect 164292 54584 164298 54596
rect 270770 54584 270776 54596
rect 164292 54556 270776 54584
rect 164292 54544 164298 54556
rect 270770 54544 270776 54556
rect 270828 54544 270834 54596
rect 313734 54544 313740 54596
rect 313792 54584 313798 54596
rect 422294 54584 422300 54596
rect 313792 54556 422300 54584
rect 313792 54544 313798 54556
rect 422294 54544 422300 54556
rect 422352 54544 422358 54596
rect 22094 54476 22100 54528
rect 22152 54516 22158 54528
rect 247402 54516 247408 54528
rect 22152 54488 247408 54516
rect 22152 54476 22158 54488
rect 247402 54476 247408 54488
rect 247460 54476 247466 54528
rect 297174 54476 297180 54528
rect 297232 54516 297238 54528
rect 322934 54516 322940 54528
rect 297232 54488 322940 54516
rect 297232 54476 297238 54488
rect 322934 54476 322940 54488
rect 322992 54476 322998 54528
rect 323670 54476 323676 54528
rect 323728 54516 323734 54528
rect 481634 54516 481640 54528
rect 323728 54488 481640 54516
rect 323728 54476 323734 54488
rect 481634 54476 481640 54488
rect 481692 54476 481698 54528
rect 166994 53116 167000 53168
rect 167052 53156 167058 53168
rect 271230 53156 271236 53168
rect 167052 53128 271236 53156
rect 167052 53116 167058 53128
rect 271230 53116 271236 53128
rect 271288 53116 271294 53168
rect 310514 53116 310520 53168
rect 310572 53156 310578 53168
rect 401686 53156 401692 53168
rect 310572 53128 401692 53156
rect 310572 53116 310578 53128
rect 401686 53116 401692 53128
rect 401744 53116 401750 53168
rect 70486 53048 70492 53100
rect 70544 53088 70550 53100
rect 255498 53088 255504 53100
rect 70544 53060 255504 53088
rect 70544 53048 70550 53060
rect 255498 53048 255504 53060
rect 255556 53048 255562 53100
rect 324314 53048 324320 53100
rect 324372 53088 324378 53100
rect 484486 53088 484492 53100
rect 324372 53060 484492 53088
rect 324372 53048 324378 53060
rect 484486 53048 484492 53060
rect 484544 53048 484550 53100
rect 175366 51756 175372 51808
rect 175424 51796 175430 51808
rect 272610 51796 272616 51808
rect 175424 51768 272616 51796
rect 175424 51756 175430 51768
rect 272610 51756 272616 51768
rect 272668 51756 272674 51808
rect 309870 51756 309876 51808
rect 309928 51796 309934 51808
rect 398834 51796 398840 51808
rect 309928 51768 398840 51796
rect 309928 51756 309934 51768
rect 398834 51756 398840 51768
rect 398892 51756 398898 51808
rect 67634 51688 67640 51740
rect 67692 51728 67698 51740
rect 254670 51728 254676 51740
rect 67692 51700 254676 51728
rect 67692 51688 67698 51700
rect 254670 51688 254676 51700
rect 254728 51688 254734 51740
rect 338850 51688 338856 51740
rect 338908 51728 338914 51740
rect 470594 51728 470600 51740
rect 338908 51700 470600 51728
rect 338908 51688 338914 51700
rect 470594 51688 470600 51700
rect 470652 51688 470658 51740
rect 178034 50396 178040 50448
rect 178092 50436 178098 50448
rect 273070 50436 273076 50448
rect 178092 50408 273076 50436
rect 178092 50396 178098 50408
rect 273070 50396 273076 50408
rect 273128 50396 273134 50448
rect 325326 50396 325332 50448
rect 325384 50436 325390 50448
rect 491294 50436 491300 50448
rect 325384 50408 491300 50436
rect 325384 50396 325390 50408
rect 491294 50396 491300 50408
rect 491352 50396 491358 50448
rect 74534 50328 74540 50380
rect 74592 50368 74598 50380
rect 255866 50368 255872 50380
rect 74592 50340 255872 50368
rect 74592 50328 74598 50340
rect 255866 50328 255872 50340
rect 255924 50328 255930 50380
rect 326062 50328 326068 50380
rect 326120 50368 326126 50380
rect 495526 50368 495532 50380
rect 326120 50340 495532 50368
rect 326120 50328 326126 50340
rect 495526 50328 495532 50340
rect 495584 50328 495590 50380
rect 3234 49648 3240 49700
rect 3292 49688 3298 49700
rect 229922 49688 229928 49700
rect 3292 49660 229928 49688
rect 3292 49648 3298 49660
rect 229922 49648 229928 49660
rect 229980 49648 229986 49700
rect 354214 49648 354220 49700
rect 354272 49688 354278 49700
rect 580166 49688 580172 49700
rect 354272 49660 580172 49688
rect 354272 49648 354278 49660
rect 580166 49648 580172 49660
rect 580224 49648 580230 49700
rect 227714 49036 227720 49088
rect 227772 49076 227778 49088
rect 281350 49076 281356 49088
rect 227772 49048 281356 49076
rect 227772 49036 227778 49048
rect 281350 49036 281356 49048
rect 281408 49036 281414 49088
rect 306006 49036 306012 49088
rect 306064 49076 306070 49088
rect 375374 49076 375380 49088
rect 306064 49048 375380 49076
rect 306064 49036 306070 49048
rect 375374 49036 375380 49048
rect 375432 49036 375438 49088
rect 131114 48968 131120 49020
rect 131172 49008 131178 49020
rect 265250 49008 265256 49020
rect 131172 48980 265256 49008
rect 131172 48968 131178 48980
rect 265250 48968 265256 48980
rect 265308 48968 265314 49020
rect 311710 48968 311716 49020
rect 311768 49008 311774 49020
rect 409874 49008 409880 49020
rect 311768 48980 409880 49008
rect 311768 48968 311774 48980
rect 409874 48968 409880 48980
rect 409932 48968 409938 49020
rect 180886 47608 180892 47660
rect 180944 47648 180950 47660
rect 273714 47648 273720 47660
rect 180944 47620 273720 47648
rect 180944 47608 180950 47620
rect 273714 47608 273720 47620
rect 273772 47608 273778 47660
rect 326430 47608 326436 47660
rect 326488 47648 326494 47660
rect 498194 47648 498200 47660
rect 326488 47620 498200 47648
rect 326488 47608 326494 47620
rect 498194 47608 498200 47620
rect 498252 47608 498258 47660
rect 93854 47540 93860 47592
rect 93912 47580 93918 47592
rect 259086 47580 259092 47592
rect 93912 47552 259092 47580
rect 93912 47540 93918 47552
rect 259086 47540 259092 47552
rect 259144 47540 259150 47592
rect 328822 47540 328828 47592
rect 328880 47580 328886 47592
rect 511994 47580 512000 47592
rect 328880 47552 512000 47580
rect 328880 47540 328886 47552
rect 511994 47540 512000 47552
rect 512052 47540 512058 47592
rect 184934 46248 184940 46300
rect 184992 46288 184998 46300
rect 274174 46288 274180 46300
rect 184992 46260 274180 46288
rect 184992 46248 184998 46260
rect 274174 46248 274180 46260
rect 274232 46248 274238 46300
rect 327074 46248 327080 46300
rect 327132 46288 327138 46300
rect 500954 46288 500960 46300
rect 327132 46260 500960 46288
rect 327132 46248 327138 46260
rect 500954 46248 500960 46260
rect 501012 46248 501018 46300
rect 31754 46180 31760 46232
rect 31812 46220 31818 46232
rect 248598 46220 248604 46232
rect 31812 46192 248604 46220
rect 31812 46180 31818 46192
rect 248598 46180 248604 46192
rect 248656 46180 248662 46232
rect 298462 46180 298468 46232
rect 298520 46220 298526 46232
rect 329834 46220 329840 46232
rect 298520 46192 329840 46220
rect 298520 46180 298526 46192
rect 329834 46180 329840 46192
rect 329892 46180 329898 46232
rect 329926 46180 329932 46232
rect 329984 46220 329990 46232
rect 518894 46220 518900 46232
rect 329984 46192 518900 46220
rect 329984 46180 329990 46192
rect 518894 46180 518900 46192
rect 518952 46180 518958 46232
rect 191926 44888 191932 44940
rect 191984 44928 191990 44940
rect 275094 44928 275100 44940
rect 191984 44900 275100 44928
rect 191984 44888 191990 44900
rect 275094 44888 275100 44900
rect 275152 44888 275158 44940
rect 328086 44888 328092 44940
rect 328144 44928 328150 44940
rect 507854 44928 507860 44940
rect 328144 44900 507860 44928
rect 328144 44888 328150 44900
rect 507854 44888 507860 44900
rect 507912 44888 507918 44940
rect 107654 44820 107660 44872
rect 107712 44860 107718 44872
rect 260926 44860 260932 44872
rect 107712 44832 260932 44860
rect 107712 44820 107718 44832
rect 260926 44820 260932 44832
rect 260984 44820 260990 44872
rect 297910 44820 297916 44872
rect 297968 44860 297974 44872
rect 327074 44860 327080 44872
rect 297968 44832 327080 44860
rect 297968 44820 297974 44832
rect 327074 44820 327080 44832
rect 327132 44820 327138 44872
rect 333790 44820 333796 44872
rect 333848 44860 333854 44872
rect 542354 44860 542360 44872
rect 333848 44832 542360 44860
rect 333848 44820 333854 44832
rect 542354 44820 542360 44832
rect 542412 44820 542418 44872
rect 142246 43460 142252 43512
rect 142304 43500 142310 43512
rect 266998 43500 267004 43512
rect 142304 43472 267004 43500
rect 142304 43460 142310 43472
rect 266998 43460 267004 43472
rect 267056 43460 267062 43512
rect 328638 43460 328644 43512
rect 328696 43500 328702 43512
rect 512086 43500 512092 43512
rect 328696 43472 512092 43500
rect 328696 43460 328702 43472
rect 512086 43460 512092 43472
rect 512144 43460 512150 43512
rect 120166 43392 120172 43444
rect 120224 43432 120230 43444
rect 263778 43432 263784 43444
rect 120224 43404 263784 43432
rect 120224 43392 120230 43404
rect 263778 43392 263784 43404
rect 263836 43392 263842 43444
rect 335446 43392 335452 43444
rect 335504 43432 335510 43444
rect 552014 43432 552020 43444
rect 335504 43404 552020 43432
rect 335504 43392 335510 43404
rect 552014 43392 552020 43404
rect 552072 43392 552078 43444
rect 204254 42100 204260 42152
rect 204312 42140 204318 42152
rect 276658 42140 276664 42152
rect 204312 42112 276664 42140
rect 204312 42100 204318 42112
rect 276658 42100 276664 42112
rect 276716 42100 276722 42152
rect 329190 42100 329196 42152
rect 329248 42140 329254 42152
rect 514754 42140 514760 42152
rect 329248 42112 514760 42140
rect 329248 42100 329254 42112
rect 514754 42100 514760 42112
rect 514812 42100 514818 42152
rect 117314 42032 117320 42084
rect 117372 42072 117378 42084
rect 262950 42072 262956 42084
rect 117372 42044 262956 42072
rect 117372 42032 117378 42044
rect 262950 42032 262956 42044
rect 263008 42032 263014 42084
rect 335998 42032 336004 42084
rect 336056 42072 336062 42084
rect 556246 42072 556252 42084
rect 336056 42044 556252 42072
rect 336056 42032 336062 42044
rect 556246 42032 556252 42044
rect 556304 42032 556310 42084
rect 301222 40808 301228 40860
rect 301280 40848 301286 40860
rect 346486 40848 346492 40860
rect 301280 40820 346492 40848
rect 301280 40808 301286 40820
rect 346486 40808 346492 40820
rect 346544 40808 346550 40860
rect 211154 40740 211160 40792
rect 211212 40780 211218 40792
rect 278590 40780 278596 40792
rect 211212 40752 278596 40780
rect 211212 40740 211218 40752
rect 278590 40740 278596 40752
rect 278648 40740 278654 40792
rect 311158 40740 311164 40792
rect 311216 40780 311222 40792
rect 407206 40780 407212 40792
rect 311216 40752 407212 40780
rect 311216 40740 311222 40752
rect 407206 40740 407212 40752
rect 407264 40740 407270 40792
rect 110414 40672 110420 40724
rect 110472 40712 110478 40724
rect 261846 40712 261852 40724
rect 110472 40684 261852 40712
rect 110472 40672 110478 40684
rect 261846 40672 261852 40684
rect 261904 40672 261910 40724
rect 331398 40672 331404 40724
rect 331456 40712 331462 40724
rect 528554 40712 528560 40724
rect 331456 40684 528560 40712
rect 331456 40672 331462 40684
rect 528554 40672 528560 40684
rect 528612 40672 528618 40724
rect 303430 39448 303436 39500
rect 303488 39488 303494 39500
rect 360194 39488 360200 39500
rect 303488 39460 360200 39488
rect 303488 39448 303494 39460
rect 360194 39448 360200 39460
rect 360252 39448 360258 39500
rect 218054 39380 218060 39432
rect 218112 39420 218118 39432
rect 279694 39420 279700 39432
rect 218112 39392 279700 39420
rect 218112 39380 218118 39392
rect 279694 39380 279700 39392
rect 279752 39380 279758 39432
rect 312814 39380 312820 39432
rect 312872 39420 312878 39432
rect 416774 39420 416780 39432
rect 312872 39392 416780 39420
rect 312872 39380 312878 39392
rect 416774 39380 416780 39392
rect 416832 39380 416838 39432
rect 84194 39312 84200 39364
rect 84252 39352 84258 39364
rect 257522 39352 257528 39364
rect 84252 39324 257528 39352
rect 84252 39312 84258 39324
rect 257522 39312 257528 39324
rect 257580 39312 257586 39364
rect 331950 39312 331956 39364
rect 332008 39352 332014 39364
rect 531314 39352 531320 39364
rect 332008 39324 531320 39352
rect 332008 39312 332014 39324
rect 531314 39312 531320 39324
rect 531372 39312 531378 39364
rect 230566 37952 230572 38004
rect 230624 37992 230630 38004
rect 281902 37992 281908 38004
rect 230624 37964 281908 37992
rect 230624 37952 230630 37964
rect 281902 37952 281908 37964
rect 281960 37952 281966 38004
rect 304534 37952 304540 38004
rect 304592 37992 304598 38004
rect 367094 37992 367100 38004
rect 304592 37964 367100 37992
rect 304592 37952 304598 37964
rect 367094 37952 367100 37964
rect 367152 37952 367158 38004
rect 38654 37884 38660 37936
rect 38712 37924 38718 37936
rect 246298 37924 246304 37936
rect 38712 37896 246304 37924
rect 38712 37884 38718 37896
rect 246298 37884 246304 37896
rect 246356 37884 246362 37936
rect 333606 37884 333612 37936
rect 333664 37924 333670 37936
rect 540974 37924 540980 37936
rect 333664 37896 540980 37924
rect 333664 37884 333670 37896
rect 540974 37884 540980 37896
rect 541032 37884 541038 37936
rect 144914 36592 144920 36644
rect 144972 36632 144978 36644
rect 267550 36632 267556 36644
rect 144972 36604 267556 36632
rect 144972 36592 144978 36604
rect 267550 36592 267556 36604
rect 267608 36592 267614 36644
rect 305086 36592 305092 36644
rect 305144 36632 305150 36644
rect 369854 36632 369860 36644
rect 305144 36604 369860 36632
rect 305144 36592 305150 36604
rect 369854 36592 369860 36604
rect 369912 36592 369918 36644
rect 44174 36524 44180 36576
rect 44232 36564 44238 36576
rect 250806 36564 250812 36576
rect 44232 36536 250812 36564
rect 44232 36524 44238 36536
rect 250806 36524 250812 36536
rect 250864 36524 250870 36576
rect 334158 36524 334164 36576
rect 334216 36564 334222 36576
rect 545206 36564 545212 36576
rect 334216 36536 545212 36564
rect 334216 36524 334222 36536
rect 545206 36524 545212 36536
rect 545264 36524 545270 36576
rect 3326 35844 3332 35896
rect 3384 35884 3390 35896
rect 229830 35884 229836 35896
rect 3384 35856 229836 35884
rect 3384 35844 3390 35856
rect 229830 35844 229836 35856
rect 229888 35844 229894 35896
rect 354122 35844 354128 35896
rect 354180 35884 354186 35896
rect 580166 35884 580172 35896
rect 354180 35856 580172 35884
rect 354180 35844 354186 35856
rect 580166 35844 580172 35856
rect 580224 35844 580230 35896
rect 299014 35232 299020 35284
rect 299072 35272 299078 35284
rect 333974 35272 333980 35284
rect 299072 35244 333980 35272
rect 299072 35232 299078 35244
rect 333974 35232 333980 35244
rect 334032 35232 334038 35284
rect 133874 35164 133880 35216
rect 133932 35204 133938 35216
rect 265802 35204 265808 35216
rect 133932 35176 265808 35204
rect 133932 35164 133938 35176
rect 265802 35164 265808 35176
rect 265860 35164 265866 35216
rect 306190 35164 306196 35216
rect 306248 35204 306254 35216
rect 376754 35204 376760 35216
rect 306248 35176 376760 35204
rect 306248 35164 306254 35176
rect 376754 35164 376760 35176
rect 376812 35164 376818 35216
rect 302326 33872 302332 33924
rect 302384 33912 302390 33924
rect 353294 33912 353300 33924
rect 302384 33884 353300 33912
rect 302384 33872 302390 33884
rect 353294 33872 353300 33884
rect 353352 33872 353358 33924
rect 151814 33804 151820 33856
rect 151872 33844 151878 33856
rect 268654 33844 268660 33856
rect 151872 33816 268660 33844
rect 151872 33804 151878 33816
rect 268654 33804 268660 33816
rect 268712 33804 268718 33856
rect 313918 33804 313924 33856
rect 313976 33844 313982 33856
rect 423766 33844 423772 33856
rect 313976 33816 423772 33844
rect 313976 33804 313982 33816
rect 423766 33804 423772 33816
rect 423824 33804 423830 33856
rect 48314 33736 48320 33788
rect 48372 33776 48378 33788
rect 251450 33776 251456 33788
rect 48372 33748 251456 33776
rect 48372 33736 48378 33748
rect 251450 33736 251456 33748
rect 251508 33736 251514 33788
rect 334710 33736 334716 33788
rect 334768 33776 334774 33788
rect 547874 33776 547880 33788
rect 334768 33748 547880 33776
rect 334768 33736 334774 33748
rect 547874 33736 547880 33748
rect 547932 33736 547938 33788
rect 92566 32444 92572 32496
rect 92624 32484 92630 32496
rect 258718 32484 258724 32496
rect 92624 32456 258724 32484
rect 92624 32444 92630 32456
rect 258718 32444 258724 32456
rect 258776 32444 258782 32496
rect 308398 32444 308404 32496
rect 308456 32484 308462 32496
rect 390646 32484 390652 32496
rect 308456 32456 390652 32484
rect 308456 32444 308462 32456
rect 390646 32444 390652 32456
rect 390704 32444 390710 32496
rect 34514 32376 34520 32428
rect 34572 32416 34578 32428
rect 235258 32416 235264 32428
rect 34572 32388 235264 32416
rect 34572 32376 34578 32388
rect 235258 32376 235264 32388
rect 235316 32376 235322 32428
rect 297358 32376 297364 32428
rect 297416 32416 297422 32428
rect 324314 32416 324320 32428
rect 297416 32388 324320 32416
rect 297416 32376 297422 32388
rect 324314 32376 324320 32388
rect 324372 32376 324378 32428
rect 336366 32376 336372 32428
rect 336424 32416 336430 32428
rect 557534 32416 557540 32428
rect 336424 32388 557540 32416
rect 336424 32376 336430 32388
rect 557534 32376 557540 32388
rect 557592 32376 557598 32428
rect 95234 31084 95240 31136
rect 95292 31124 95298 31136
rect 259270 31124 259276 31136
rect 95292 31096 259276 31124
rect 95292 31084 95298 31096
rect 259270 31084 259276 31096
rect 259328 31084 259334 31136
rect 311526 31084 311532 31136
rect 311584 31124 311590 31136
rect 408494 31124 408500 31136
rect 311584 31096 408500 31124
rect 311584 31084 311590 31096
rect 408494 31084 408500 31096
rect 408552 31084 408558 31136
rect 32398 31016 32404 31068
rect 32456 31056 32462 31068
rect 247862 31056 247868 31068
rect 32456 31028 247868 31056
rect 32456 31016 32462 31028
rect 247862 31016 247868 31028
rect 247920 31016 247926 31068
rect 323302 31016 323308 31068
rect 323360 31056 323366 31068
rect 478966 31056 478972 31068
rect 323360 31028 478972 31056
rect 323360 31016 323366 31028
rect 478966 31016 478972 31028
rect 479024 31016 479030 31068
rect 102134 29656 102140 29708
rect 102192 29696 102198 29708
rect 260374 29696 260380 29708
rect 102192 29668 260380 29696
rect 102192 29656 102198 29668
rect 260374 29656 260380 29668
rect 260432 29656 260438 29708
rect 312630 29656 312636 29708
rect 312688 29696 312694 29708
rect 415394 29696 415400 29708
rect 312688 29668 415400 29696
rect 312688 29656 312694 29668
rect 415394 29656 415400 29668
rect 415452 29656 415458 29708
rect 64874 29588 64880 29640
rect 64932 29628 64938 29640
rect 254118 29628 254124 29640
rect 64932 29600 254124 29628
rect 64932 29588 64938 29600
rect 254118 29588 254124 29600
rect 254176 29588 254182 29640
rect 323854 29588 323860 29640
rect 323912 29628 323918 29640
rect 483014 29628 483020 29640
rect 323912 29600 483020 29628
rect 323912 29588 323918 29600
rect 483014 29588 483020 29600
rect 483072 29588 483078 29640
rect 111794 28296 111800 28348
rect 111852 28336 111858 28348
rect 262030 28336 262036 28348
rect 111852 28308 262036 28336
rect 111852 28296 111858 28308
rect 262030 28296 262036 28308
rect 262088 28296 262094 28348
rect 314286 28296 314292 28348
rect 314344 28336 314350 28348
rect 425054 28336 425060 28348
rect 314344 28308 425060 28336
rect 314344 28296 314350 28308
rect 425054 28296 425060 28308
rect 425112 28296 425118 28348
rect 77294 28228 77300 28280
rect 77352 28268 77358 28280
rect 256326 28268 256332 28280
rect 77352 28240 256332 28268
rect 77352 28228 77358 28240
rect 256326 28228 256332 28240
rect 256384 28228 256390 28280
rect 324958 28228 324964 28280
rect 325016 28268 325022 28280
rect 490006 28268 490012 28280
rect 325016 28240 490012 28268
rect 325016 28228 325022 28240
rect 490006 28228 490012 28240
rect 490064 28228 490070 28280
rect 114646 26936 114652 26988
rect 114704 26976 114710 26988
rect 262674 26976 262680 26988
rect 114704 26948 262680 26976
rect 114704 26936 114710 26948
rect 262674 26936 262680 26948
rect 262732 26936 262738 26988
rect 314838 26936 314844 26988
rect 314896 26976 314902 26988
rect 429286 26976 429292 26988
rect 314896 26948 429292 26976
rect 314896 26936 314902 26948
rect 429286 26936 429292 26948
rect 429344 26936 429350 26988
rect 81526 26868 81532 26920
rect 81584 26908 81590 26920
rect 257154 26908 257160 26920
rect 81584 26880 257160 26908
rect 81584 26868 81590 26880
rect 257154 26868 257160 26880
rect 257212 26868 257218 26920
rect 325510 26868 325516 26920
rect 325568 26908 325574 26920
rect 492674 26908 492680 26920
rect 325568 26880 492680 26908
rect 325568 26868 325574 26880
rect 492674 26868 492680 26880
rect 492732 26868 492738 26920
rect 125686 25576 125692 25628
rect 125744 25616 125750 25628
rect 264330 25616 264336 25628
rect 125744 25588 264336 25616
rect 125744 25576 125750 25588
rect 264330 25576 264336 25588
rect 264388 25576 264394 25628
rect 315390 25576 315396 25628
rect 315448 25616 315454 25628
rect 431954 25616 431960 25628
rect 315448 25588 431960 25616
rect 315448 25576 315454 25588
rect 431954 25576 431960 25588
rect 432012 25576 432018 25628
rect 98086 25508 98092 25560
rect 98144 25548 98150 25560
rect 259546 25548 259552 25560
rect 98144 25520 259552 25548
rect 98144 25508 98150 25520
rect 259546 25508 259552 25520
rect 259604 25508 259610 25560
rect 326614 25508 326620 25560
rect 326672 25548 326678 25560
rect 499574 25548 499580 25560
rect 326672 25520 499580 25548
rect 326672 25508 326678 25520
rect 499574 25508 499580 25520
rect 499632 25508 499638 25560
rect 118694 24148 118700 24200
rect 118752 24188 118758 24200
rect 263134 24188 263140 24200
rect 118752 24160 263140 24188
rect 118752 24148 118758 24160
rect 263134 24148 263140 24160
rect 263192 24148 263198 24200
rect 317598 24148 317604 24200
rect 317656 24188 317662 24200
rect 445846 24188 445852 24200
rect 317656 24160 445852 24188
rect 317656 24148 317662 24160
rect 445846 24148 445852 24160
rect 445904 24148 445910 24200
rect 87046 24080 87052 24132
rect 87104 24120 87110 24132
rect 257338 24120 257344 24132
rect 87104 24092 257344 24120
rect 87104 24080 87110 24092
rect 257338 24080 257344 24092
rect 257396 24080 257402 24132
rect 327718 24080 327724 24132
rect 327776 24120 327782 24132
rect 506566 24120 506572 24132
rect 327776 24092 506572 24120
rect 327776 24080 327782 24092
rect 506566 24080 506572 24092
rect 506624 24080 506630 24132
rect 354030 23400 354036 23452
rect 354088 23440 354094 23452
rect 580166 23440 580172 23452
rect 354088 23412 580172 23440
rect 354088 23400 354094 23412
rect 580166 23400 580172 23412
rect 580224 23400 580230 23452
rect 168374 22788 168380 22840
rect 168432 22828 168438 22840
rect 271414 22828 271420 22840
rect 168432 22800 271420 22828
rect 168432 22788 168438 22800
rect 271414 22788 271420 22800
rect 271472 22788 271478 22840
rect 299566 22788 299572 22840
rect 299624 22828 299630 22840
rect 336826 22828 336832 22840
rect 299624 22800 336832 22828
rect 299624 22788 299630 22800
rect 336826 22788 336832 22800
rect 336884 22788 336890 22840
rect 60734 22720 60740 22772
rect 60792 22760 60798 22772
rect 253566 22760 253572 22772
rect 60792 22732 253572 22760
rect 60792 22720 60798 22732
rect 253566 22720 253572 22732
rect 253624 22720 253630 22772
rect 307294 22720 307300 22772
rect 307352 22760 307358 22772
rect 383654 22760 383660 22772
rect 307352 22732 383660 22760
rect 307352 22720 307358 22732
rect 383654 22720 383660 22732
rect 383712 22720 383718 22772
rect 164326 21428 164332 21480
rect 164384 21468 164390 21480
rect 270954 21468 270960 21480
rect 164384 21440 270960 21468
rect 164384 21428 164390 21440
rect 270954 21428 270960 21440
rect 271012 21428 271018 21480
rect 318150 21428 318156 21480
rect 318208 21468 318214 21480
rect 448514 21468 448520 21480
rect 318208 21440 448520 21468
rect 318208 21428 318214 21440
rect 448514 21428 448520 21440
rect 448572 21428 448578 21480
rect 27614 21360 27620 21412
rect 27672 21400 27678 21412
rect 248046 21400 248052 21412
rect 27672 21372 248052 21400
rect 27672 21360 27678 21372
rect 248046 21360 248052 21372
rect 248104 21360 248110 21412
rect 328270 21360 328276 21412
rect 328328 21400 328334 21412
rect 509234 21400 509240 21412
rect 328328 21372 509240 21400
rect 328328 21360 328334 21372
rect 509234 21360 509240 21372
rect 509292 21360 509298 21412
rect 154574 20000 154580 20052
rect 154632 20040 154638 20052
rect 269206 20040 269212 20052
rect 154632 20012 269212 20040
rect 154632 20000 154638 20012
rect 269206 20000 269212 20012
rect 269264 20000 269270 20052
rect 319806 20000 319812 20052
rect 319864 20040 319870 20052
rect 458174 20040 458180 20052
rect 319864 20012 458180 20040
rect 319864 20000 319870 20012
rect 458174 20000 458180 20012
rect 458232 20000 458238 20052
rect 71774 19932 71780 19984
rect 71832 19972 71838 19984
rect 255406 19972 255412 19984
rect 71832 19944 255412 19972
rect 71832 19932 71838 19944
rect 255406 19932 255412 19944
rect 255464 19932 255470 19984
rect 330478 19932 330484 19984
rect 330536 19972 330542 19984
rect 523034 19972 523040 19984
rect 330536 19944 523040 19972
rect 330536 19932 330542 19944
rect 523034 19932 523040 19944
rect 523092 19932 523098 19984
rect 147766 18640 147772 18692
rect 147824 18680 147830 18692
rect 268286 18680 268292 18692
rect 147824 18652 268292 18680
rect 147824 18640 147830 18652
rect 268286 18640 268292 18652
rect 268344 18640 268350 18692
rect 320910 18640 320916 18692
rect 320968 18680 320974 18692
rect 465074 18680 465080 18692
rect 320968 18652 465080 18680
rect 320968 18640 320974 18652
rect 465074 18640 465080 18652
rect 465132 18640 465138 18692
rect 76006 18572 76012 18624
rect 76064 18612 76070 18624
rect 256050 18612 256056 18624
rect 76064 18584 256056 18612
rect 76064 18572 76070 18584
rect 256050 18572 256056 18584
rect 256108 18572 256114 18624
rect 331582 18572 331588 18624
rect 331640 18612 331646 18624
rect 528646 18612 528652 18624
rect 331640 18584 528652 18612
rect 331640 18572 331646 18584
rect 528646 18572 528652 18584
rect 528704 18572 528710 18624
rect 244274 17348 244280 17400
rect 244332 17388 244338 17400
rect 284110 17388 284116 17400
rect 244332 17360 284116 17388
rect 244332 17348 244338 17360
rect 284110 17348 284116 17360
rect 284168 17348 284174 17400
rect 109126 17280 109132 17332
rect 109184 17320 109190 17332
rect 261570 17320 261576 17332
rect 109184 17292 261576 17320
rect 109184 17280 109190 17292
rect 261570 17280 261576 17292
rect 261628 17280 261634 17332
rect 321646 17280 321652 17332
rect 321704 17320 321710 17332
rect 469214 17320 469220 17332
rect 321704 17292 469220 17320
rect 321704 17280 321710 17292
rect 469214 17280 469220 17292
rect 469272 17280 469278 17332
rect 73154 17212 73160 17264
rect 73212 17252 73218 17264
rect 244918 17252 244924 17264
rect 73212 17224 244924 17252
rect 73212 17212 73218 17224
rect 244918 17212 244924 17224
rect 244976 17212 244982 17264
rect 333238 17212 333244 17264
rect 333296 17252 333302 17264
rect 539686 17252 539692 17264
rect 333296 17224 539692 17252
rect 333296 17212 333302 17224
rect 539686 17212 539692 17224
rect 539744 17212 539750 17264
rect 241698 15920 241704 15972
rect 241756 15960 241762 15972
rect 283374 15960 283380 15972
rect 241756 15932 283380 15960
rect 241756 15920 241762 15932
rect 283374 15920 283380 15932
rect 283432 15920 283438 15972
rect 322198 15920 322204 15972
rect 322256 15960 322262 15972
rect 473538 15960 473544 15972
rect 322256 15932 473544 15960
rect 322256 15920 322262 15932
rect 473538 15920 473544 15932
rect 473596 15920 473602 15972
rect 101490 15852 101496 15904
rect 101548 15892 101554 15904
rect 260190 15892 260196 15904
rect 101548 15864 260196 15892
rect 101548 15852 101554 15864
rect 260190 15852 260196 15864
rect 260248 15852 260254 15904
rect 334894 15852 334900 15904
rect 334952 15892 334958 15904
rect 549714 15892 549720 15904
rect 334952 15864 549720 15892
rect 334952 15852 334958 15864
rect 549714 15852 549720 15864
rect 549772 15852 549778 15904
rect 208578 14492 208584 14544
rect 208636 14532 208642 14544
rect 277854 14532 277860 14544
rect 208636 14504 277860 14532
rect 208636 14492 208642 14504
rect 277854 14492 277860 14504
rect 277912 14492 277918 14544
rect 325050 14492 325056 14544
rect 325108 14532 325114 14544
rect 451366 14532 451372 14544
rect 325108 14504 451372 14532
rect 325108 14492 325114 14504
rect 451366 14492 451372 14504
rect 451424 14492 451430 14544
rect 124674 14424 124680 14476
rect 124732 14464 124738 14476
rect 263686 14464 263692 14476
rect 124732 14436 263692 14464
rect 124732 14424 124738 14436
rect 263686 14424 263692 14436
rect 263744 14424 263750 14476
rect 295150 14424 295156 14476
rect 295208 14464 295214 14476
rect 311250 14464 311256 14476
rect 295208 14436 311256 14464
rect 295208 14424 295214 14436
rect 311250 14424 311256 14436
rect 311308 14424 311314 14476
rect 329374 14424 329380 14476
rect 329432 14464 329438 14476
rect 516594 14464 516600 14476
rect 329432 14436 516600 14464
rect 329432 14424 329438 14436
rect 516594 14424 516600 14436
rect 516652 14424 516658 14476
rect 195330 13132 195336 13184
rect 195388 13172 195394 13184
rect 275830 13172 275836 13184
rect 195388 13144 275836 13172
rect 195388 13132 195394 13144
rect 275830 13132 275836 13144
rect 275888 13132 275894 13184
rect 308950 13132 308956 13184
rect 309008 13172 309014 13184
rect 394050 13172 394056 13184
rect 309008 13144 394056 13172
rect 309008 13132 309014 13144
rect 394050 13132 394056 13144
rect 394108 13132 394114 13184
rect 127986 13064 127992 13116
rect 128044 13104 128050 13116
rect 264606 13104 264612 13116
rect 128044 13076 264612 13104
rect 128044 13064 128050 13076
rect 264606 13064 264612 13076
rect 264664 13064 264670 13116
rect 298278 13064 298284 13116
rect 298336 13104 298342 13116
rect 330018 13104 330024 13116
rect 298336 13076 330024 13104
rect 298336 13064 298342 13076
rect 330018 13064 330024 13076
rect 330076 13064 330082 13116
rect 340138 13064 340144 13116
rect 340196 13104 340202 13116
rect 550726 13104 550732 13116
rect 340196 13076 550732 13104
rect 340196 13064 340202 13076
rect 550726 13064 550732 13076
rect 550784 13064 550790 13116
rect 158898 11772 158904 11824
rect 158956 11812 158962 11824
rect 269758 11812 269764 11824
rect 158956 11784 269764 11812
rect 158956 11772 158962 11784
rect 269758 11772 269764 11784
rect 269816 11772 269822 11824
rect 306742 11772 306748 11824
rect 306800 11812 306806 11824
rect 379606 11812 379612 11824
rect 306800 11784 379612 11812
rect 306800 11772 306806 11784
rect 379606 11772 379612 11784
rect 379664 11772 379670 11824
rect 69474 11704 69480 11756
rect 69532 11744 69538 11756
rect 254854 11744 254860 11756
rect 69532 11716 254860 11744
rect 69532 11704 69538 11716
rect 254854 11704 254860 11716
rect 254912 11704 254918 11756
rect 263778 11704 263784 11756
rect 263836 11744 263842 11756
rect 286318 11744 286324 11756
rect 263836 11716 286324 11744
rect 263836 11704 263842 11716
rect 286318 11704 286324 11716
rect 286376 11704 286382 11756
rect 297726 11704 297732 11756
rect 297784 11744 297790 11756
rect 326706 11744 326712 11756
rect 297784 11716 326712 11744
rect 297784 11704 297790 11716
rect 326706 11704 326712 11716
rect 326764 11704 326770 11756
rect 338758 11704 338764 11756
rect 338816 11744 338822 11756
rect 537570 11744 537576 11756
rect 338816 11716 537576 11744
rect 338816 11704 338822 11716
rect 537570 11704 537576 11716
rect 537628 11704 537634 11756
rect 300210 10956 300216 11008
rect 300268 10996 300274 11008
rect 304166 10996 304172 11008
rect 300268 10968 304172 10996
rect 300268 10956 300274 10968
rect 304166 10956 304172 10968
rect 304224 10956 304230 11008
rect 186498 10344 186504 10396
rect 186556 10384 186562 10396
rect 239398 10384 239404 10396
rect 186556 10356 239404 10384
rect 186556 10344 186562 10356
rect 239398 10344 239404 10356
rect 239456 10344 239462 10396
rect 247402 10344 247408 10396
rect 247460 10384 247466 10396
rect 284662 10384 284668 10396
rect 247460 10356 284668 10384
rect 247460 10344 247466 10356
rect 284662 10344 284668 10356
rect 284720 10344 284726 10396
rect 310054 10344 310060 10396
rect 310112 10384 310118 10396
rect 400674 10384 400680 10396
rect 310112 10356 400680 10384
rect 310112 10344 310118 10356
rect 400674 10344 400680 10356
rect 400732 10344 400738 10396
rect 51810 10276 51816 10328
rect 51868 10316 51874 10328
rect 251910 10316 251916 10328
rect 51868 10288 251916 10316
rect 51868 10276 51874 10288
rect 251910 10276 251916 10288
rect 251968 10276 251974 10328
rect 257154 10276 257160 10328
rect 257212 10316 257218 10328
rect 286134 10316 286140 10328
rect 257212 10288 286140 10316
rect 257212 10276 257218 10288
rect 286134 10276 286140 10288
rect 286192 10276 286198 10328
rect 293310 10276 293316 10328
rect 293368 10316 293374 10328
rect 300210 10316 300216 10328
rect 293368 10288 300216 10316
rect 293368 10276 293374 10288
rect 300210 10276 300216 10288
rect 300268 10276 300274 10328
rect 300670 10276 300676 10328
rect 300728 10316 300734 10328
rect 344370 10316 344376 10328
rect 300728 10288 344376 10316
rect 300728 10276 300734 10288
rect 344370 10276 344376 10288
rect 344428 10276 344434 10328
rect 347038 10276 347044 10328
rect 347096 10316 347102 10328
rect 523126 10316 523132 10328
rect 347096 10288 523132 10316
rect 347096 10276 347102 10288
rect 523126 10276 523132 10288
rect 523184 10276 523190 10328
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 229738 9636 229744 9648
rect 3476 9608 229744 9636
rect 3476 9596 3482 9608
rect 229738 9596 229744 9608
rect 229796 9596 229802 9648
rect 353938 9596 353944 9648
rect 353996 9636 354002 9648
rect 580166 9636 580172 9648
rect 353996 9608 580172 9636
rect 353996 9596 354002 9608
rect 580166 9596 580172 9608
rect 580224 9596 580230 9648
rect 229554 9528 229560 9580
rect 229612 9568 229618 9580
rect 238018 9568 238024 9580
rect 229612 9540 238024 9568
rect 229612 9528 229618 9540
rect 238018 9528 238024 9540
rect 238076 9528 238082 9580
rect 105906 9120 105912 9172
rect 105964 9160 105970 9172
rect 261478 9160 261484 9172
rect 105964 9132 261484 9160
rect 105964 9120 105970 9132
rect 261478 9120 261484 9132
rect 261536 9120 261542 9172
rect 279234 9120 279240 9172
rect 279292 9160 279298 9172
rect 289170 9160 289176 9172
rect 279292 9132 289176 9160
rect 279292 9120 279298 9132
rect 289170 9120 289176 9132
rect 289228 9120 289234 9172
rect 260466 9052 260472 9104
rect 260524 9092 260530 9104
rect 286686 9092 286692 9104
rect 260524 9064 286692 9092
rect 260524 9052 260530 9064
rect 286686 9052 286692 9064
rect 286744 9052 286750 9104
rect 247218 8984 247224 9036
rect 247276 9024 247282 9036
rect 283650 9024 283656 9036
rect 247276 8996 283656 9024
rect 247276 8984 247282 8996
rect 283650 8984 283656 8996
rect 283708 8984 283714 9036
rect 296714 8984 296720 9036
rect 296772 9024 296778 9036
rect 320082 9024 320088 9036
rect 296772 8996 320088 9024
rect 296772 8984 296778 8996
rect 320082 8984 320088 8996
rect 320140 8984 320146 9036
rect 261570 8916 261576 8968
rect 261628 8956 261634 8968
rect 286870 8956 286876 8968
rect 261628 8928 286876 8956
rect 261628 8916 261634 8928
rect 286870 8916 286876 8928
rect 286928 8916 286934 8968
rect 302878 8916 302884 8968
rect 302936 8956 302942 8968
rect 357618 8956 357624 8968
rect 302936 8928 357624 8956
rect 302936 8916 302942 8928
rect 357618 8916 357624 8928
rect 357676 8916 357682 8968
rect 251634 7692 251640 7744
rect 251692 7732 251698 7744
rect 285214 7732 285220 7744
rect 251692 7704 285220 7732
rect 251692 7692 251698 7704
rect 285214 7692 285220 7704
rect 285272 7692 285278 7744
rect 173250 7624 173256 7676
rect 173308 7664 173314 7676
rect 242158 7664 242164 7676
rect 173308 7636 242164 7664
rect 173308 7624 173314 7636
rect 242158 7624 242164 7636
rect 242216 7624 242222 7676
rect 250530 7624 250536 7676
rect 250588 7664 250594 7676
rect 285030 7664 285036 7676
rect 250588 7636 285036 7664
rect 250588 7624 250594 7636
rect 285030 7624 285036 7636
rect 285088 7624 285094 7676
rect 305638 7624 305644 7676
rect 305696 7664 305702 7676
rect 374178 7664 374184 7676
rect 305696 7636 374184 7664
rect 305696 7624 305702 7636
rect 374178 7624 374184 7636
rect 374236 7624 374242 7676
rect 66162 7556 66168 7608
rect 66220 7596 66226 7608
rect 254394 7596 254400 7608
rect 66220 7568 254400 7596
rect 66220 7556 66226 7568
rect 254394 7556 254400 7568
rect 254452 7556 254458 7608
rect 265986 7556 265992 7608
rect 266044 7596 266050 7608
rect 287146 7596 287152 7608
rect 266044 7568 287152 7596
rect 266044 7556 266050 7568
rect 287146 7556 287152 7568
rect 287204 7556 287210 7608
rect 296438 7556 296444 7608
rect 296496 7596 296502 7608
rect 318978 7596 318984 7608
rect 296496 7568 318984 7596
rect 296496 7556 296502 7568
rect 318978 7556 318984 7568
rect 319036 7556 319042 7608
rect 345658 7556 345664 7608
rect 345716 7596 345722 7608
rect 501138 7596 501144 7608
rect 345716 7568 501144 7596
rect 345716 7556 345722 7568
rect 501138 7556 501144 7568
rect 501196 7556 501202 7608
rect 275922 6876 275928 6928
rect 275980 6916 275986 6928
rect 279510 6916 279516 6928
rect 275980 6888 279516 6916
rect 275980 6876 275986 6888
rect 279510 6876 279516 6888
rect 279568 6876 279574 6928
rect 270402 6400 270408 6452
rect 270460 6440 270466 6452
rect 278038 6440 278044 6452
rect 270460 6412 278044 6440
rect 270460 6400 270466 6412
rect 278038 6400 278044 6412
rect 278096 6400 278102 6452
rect 253842 6332 253848 6384
rect 253900 6372 253906 6384
rect 275278 6372 275284 6384
rect 253900 6344 275284 6372
rect 253900 6332 253906 6344
rect 275278 6332 275284 6344
rect 275336 6332 275342 6384
rect 262674 6264 262680 6316
rect 262732 6304 262738 6316
rect 284938 6304 284944 6316
rect 262732 6276 284944 6304
rect 262732 6264 262738 6276
rect 284938 6264 284944 6276
rect 284996 6264 285002 6316
rect 304442 6264 304448 6316
rect 304500 6304 304506 6316
rect 313458 6304 313464 6316
rect 304500 6276 313464 6304
rect 304500 6264 304506 6276
rect 313458 6264 313464 6276
rect 313516 6264 313522 6316
rect 20898 6196 20904 6248
rect 20956 6236 20962 6248
rect 245746 6236 245752 6248
rect 20956 6208 245752 6236
rect 20956 6196 20962 6208
rect 245746 6196 245752 6208
rect 245804 6196 245810 6248
rect 258258 6196 258264 6248
rect 258316 6236 258322 6248
rect 286410 6236 286416 6248
rect 258316 6208 286416 6236
rect 258316 6196 258322 6208
rect 286410 6196 286416 6208
rect 286468 6196 286474 6248
rect 294598 6196 294604 6248
rect 294656 6236 294662 6248
rect 307938 6236 307944 6248
rect 294656 6208 307944 6236
rect 294656 6196 294662 6208
rect 307938 6196 307944 6208
rect 307996 6196 308002 6248
rect 342898 6196 342904 6248
rect 342956 6236 342962 6248
rect 487890 6236 487896 6248
rect 342956 6208 487896 6236
rect 342956 6196 342962 6208
rect 487890 6196 487896 6208
rect 487948 6196 487954 6248
rect 19794 6128 19800 6180
rect 19852 6168 19858 6180
rect 245654 6168 245660 6180
rect 19852 6140 245660 6168
rect 19852 6128 19858 6140
rect 245654 6128 245660 6140
rect 245712 6128 245718 6180
rect 252738 6128 252744 6180
rect 252796 6168 252802 6180
rect 285398 6168 285404 6180
rect 252796 6140 285404 6168
rect 252796 6128 252802 6140
rect 285398 6128 285404 6140
rect 285456 6128 285462 6180
rect 285858 6128 285864 6180
rect 285916 6168 285922 6180
rect 290918 6168 290924 6180
rect 285916 6140 290924 6168
rect 285916 6128 285922 6140
rect 290918 6128 290924 6140
rect 290976 6128 290982 6180
rect 295886 6128 295892 6180
rect 295944 6168 295950 6180
rect 315666 6168 315672 6180
rect 295944 6140 315672 6168
rect 295944 6128 295950 6140
rect 315666 6128 315672 6140
rect 315724 6128 315730 6180
rect 332134 6128 332140 6180
rect 332192 6168 332198 6180
rect 533154 6168 533160 6180
rect 332192 6140 533160 6168
rect 332192 6128 332198 6140
rect 533154 6128 533160 6140
rect 533212 6128 533218 6180
rect 280338 5516 280344 5568
rect 280396 5556 280402 5568
rect 289078 5556 289084 5568
rect 280396 5528 289084 5556
rect 280396 5516 280402 5528
rect 289078 5516 289084 5528
rect 289136 5516 289142 5568
rect 272610 5108 272616 5160
rect 272668 5148 272674 5160
rect 282270 5148 282276 5160
rect 272668 5120 282276 5148
rect 272668 5108 272674 5120
rect 282270 5108 282276 5120
rect 282328 5108 282334 5160
rect 269298 5040 269304 5092
rect 269356 5080 269362 5092
rect 288158 5080 288164 5092
rect 269356 5052 288164 5080
rect 269356 5040 269362 5052
rect 288158 5040 288164 5052
rect 288216 5040 288222 5092
rect 256050 4972 256056 5024
rect 256108 5012 256114 5024
rect 273898 5012 273904 5024
rect 256108 4984 273904 5012
rect 256108 4972 256114 4984
rect 273898 4972 273904 4984
rect 273956 4972 273962 5024
rect 136818 4904 136824 4956
rect 136876 4944 136882 4956
rect 136876 4916 142154 4944
rect 136876 4904 136882 4916
rect 142126 4876 142154 4916
rect 254946 4904 254952 4956
rect 255004 4944 255010 4956
rect 283558 4944 283564 4956
rect 255004 4916 283564 4944
rect 255004 4904 255010 4916
rect 283558 4904 283564 4916
rect 283616 4904 283622 4956
rect 293678 4904 293684 4956
rect 293736 4944 293742 4956
rect 302418 4944 302424 4956
rect 293736 4916 302424 4944
rect 293736 4904 293742 4916
rect 302418 4904 302424 4916
rect 302476 4904 302482 4956
rect 243538 4876 243544 4888
rect 142126 4848 243544 4876
rect 243538 4836 243544 4848
rect 243596 4836 243602 4888
rect 249426 4836 249432 4888
rect 249484 4876 249490 4888
rect 282178 4876 282184 4888
rect 249484 4848 282184 4876
rect 249484 4836 249490 4848
rect 282178 4836 282184 4848
rect 282236 4836 282242 4888
rect 295334 4836 295340 4888
rect 295392 4876 295398 4888
rect 312354 4876 312360 4888
rect 295392 4848 312360 4876
rect 295392 4836 295398 4848
rect 312354 4836 312360 4848
rect 312412 4836 312418 4888
rect 341518 4836 341524 4888
rect 341576 4876 341582 4888
rect 474642 4876 474648 4888
rect 341576 4848 474648 4876
rect 341576 4836 341582 4848
rect 474642 4836 474648 4848
rect 474700 4836 474706 4888
rect 475378 4836 475384 4888
rect 475436 4876 475442 4888
rect 497826 4876 497832 4888
rect 475436 4848 497832 4876
rect 475436 4836 475442 4848
rect 497826 4836 497832 4848
rect 497884 4836 497890 4888
rect 86034 4768 86040 4820
rect 86092 4808 86098 4820
rect 257614 4808 257620 4820
rect 86092 4780 257620 4808
rect 86092 4768 86098 4780
rect 257614 4768 257620 4780
rect 257672 4768 257678 4820
rect 259362 4768 259368 4820
rect 259420 4808 259426 4820
rect 279418 4808 279424 4820
rect 259420 4780 279424 4808
rect 259420 4768 259426 4780
rect 279418 4768 279424 4780
rect 279476 4768 279482 4820
rect 296070 4768 296076 4820
rect 296128 4808 296134 4820
rect 316770 4808 316776 4820
rect 296128 4780 316776 4808
rect 296128 4768 296134 4780
rect 316770 4768 316776 4780
rect 316828 4768 316834 4820
rect 323762 4768 323768 4820
rect 323820 4808 323826 4820
rect 335538 4808 335544 4820
rect 323820 4780 335544 4808
rect 323820 4768 323826 4780
rect 335538 4768 335544 4780
rect 335596 4768 335602 4820
rect 336550 4768 336556 4820
rect 336608 4808 336614 4820
rect 559650 4808 559656 4820
rect 336608 4780 559656 4808
rect 336608 4768 336614 4780
rect 559650 4768 559656 4780
rect 559708 4768 559714 4820
rect 301682 4496 301688 4548
rect 301740 4536 301746 4548
rect 309042 4536 309048 4548
rect 301740 4508 309048 4536
rect 301740 4496 301746 4508
rect 309042 4496 309048 4508
rect 309100 4496 309106 4548
rect 282546 4428 282552 4480
rect 282604 4468 282610 4480
rect 287698 4468 287704 4480
rect 282604 4440 287704 4468
rect 282604 4428 282610 4440
rect 287698 4428 287704 4440
rect 287756 4428 287762 4480
rect 293126 4360 293132 4412
rect 293184 4400 293190 4412
rect 299106 4400 299112 4412
rect 293184 4372 299112 4400
rect 293184 4360 293190 4372
rect 299106 4360 299112 4372
rect 299164 4360 299170 4412
rect 70486 4156 70492 4208
rect 70544 4196 70550 4208
rect 71682 4196 71688 4208
rect 70544 4168 71688 4196
rect 70544 4156 70550 4168
rect 71682 4156 71688 4168
rect 71740 4156 71746 4208
rect 87046 4156 87052 4208
rect 87104 4196 87110 4208
rect 88242 4196 88248 4208
rect 87104 4168 88248 4196
rect 87104 4156 87110 4168
rect 88242 4156 88248 4168
rect 88300 4156 88306 4208
rect 114646 4156 114652 4208
rect 114704 4196 114710 4208
rect 115842 4196 115848 4208
rect 114704 4168 115848 4196
rect 114704 4156 114710 4168
rect 115842 4156 115848 4168
rect 115900 4156 115906 4208
rect 120166 4156 120172 4208
rect 120224 4196 120230 4208
rect 121362 4196 121368 4208
rect 120224 4168 121368 4196
rect 120224 4156 120230 4168
rect 121362 4156 121368 4168
rect 121420 4156 121426 4208
rect 147766 4156 147772 4208
rect 147824 4196 147830 4208
rect 148962 4196 148968 4208
rect 147824 4168 148968 4196
rect 147824 4156 147830 4168
rect 148962 4156 148968 4168
rect 149020 4156 149026 4208
rect 153286 4156 153292 4208
rect 153344 4196 153350 4208
rect 154482 4196 154488 4208
rect 153344 4168 154488 4196
rect 153344 4156 153350 4168
rect 154482 4156 154488 4168
rect 154540 4156 154546 4208
rect 164326 4156 164332 4208
rect 164384 4196 164390 4208
rect 165522 4196 165528 4208
rect 164384 4168 165528 4196
rect 164384 4156 164390 4168
rect 165522 4156 165528 4168
rect 165580 4156 165586 4208
rect 169846 4156 169852 4208
rect 169904 4196 169910 4208
rect 171042 4196 171048 4208
rect 169904 4168 171048 4196
rect 169904 4156 169910 4168
rect 171042 4156 171048 4168
rect 171100 4156 171106 4208
rect 180886 4156 180892 4208
rect 180944 4196 180950 4208
rect 182082 4196 182088 4208
rect 180944 4168 182088 4196
rect 180944 4156 180950 4168
rect 182082 4156 182088 4168
rect 182140 4156 182146 4208
rect 197446 4156 197452 4208
rect 197504 4196 197510 4208
rect 198642 4196 198648 4208
rect 197504 4168 198648 4196
rect 197504 4156 197510 4168
rect 198642 4156 198648 4168
rect 198700 4156 198706 4208
rect 202966 4156 202972 4208
rect 203024 4196 203030 4208
rect 204162 4196 204168 4208
rect 203024 4168 204168 4196
rect 203024 4156 203030 4168
rect 204162 4156 204168 4168
rect 204220 4156 204226 4208
rect 214006 4156 214012 4208
rect 214064 4196 214070 4208
rect 215202 4196 215208 4208
rect 214064 4168 215208 4196
rect 214064 4156 214070 4168
rect 215202 4156 215208 4168
rect 215260 4156 215266 4208
rect 230566 4156 230572 4208
rect 230624 4196 230630 4208
rect 231762 4196 231768 4208
rect 230624 4168 231768 4196
rect 230624 4156 230630 4168
rect 231762 4156 231768 4168
rect 231820 4156 231826 4208
rect 236086 4156 236092 4208
rect 236144 4196 236150 4208
rect 237282 4196 237288 4208
rect 236144 4168 237288 4196
rect 236144 4156 236150 4168
rect 237282 4156 237288 4168
rect 237340 4156 237346 4208
rect 301498 4156 301504 4208
rect 301556 4196 301562 4208
rect 303522 4196 303528 4208
rect 301556 4168 303528 4196
rect 301556 4156 301562 4168
rect 303522 4156 303528 4168
rect 303580 4156 303586 4208
rect 304258 4156 304264 4208
rect 304316 4196 304322 4208
rect 305730 4196 305736 4208
rect 304316 4168 305736 4196
rect 304316 4156 304322 4168
rect 305730 4156 305736 4168
rect 305788 4156 305794 4208
rect 320818 4156 320824 4208
rect 320876 4196 320882 4208
rect 322290 4196 322296 4208
rect 320876 4168 322296 4196
rect 320876 4156 320882 4168
rect 322290 4156 322296 4168
rect 322348 4156 322354 4208
rect 323578 4156 323584 4208
rect 323636 4196 323642 4208
rect 325602 4196 325608 4208
rect 323636 4168 325608 4196
rect 323636 4156 323642 4168
rect 325602 4156 325608 4168
rect 325660 4156 325666 4208
rect 346486 4156 346492 4208
rect 346544 4196 346550 4208
rect 347682 4196 347688 4208
rect 346544 4168 347688 4196
rect 346544 4156 346550 4168
rect 347682 4156 347688 4168
rect 347740 4156 347746 4208
rect 352006 4156 352012 4208
rect 352064 4196 352070 4208
rect 353202 4196 353208 4208
rect 352064 4168 353208 4196
rect 352064 4156 352070 4168
rect 353202 4156 353208 4168
rect 353260 4156 353266 4208
rect 363046 4156 363052 4208
rect 363104 4196 363110 4208
rect 364242 4196 364248 4208
rect 363104 4168 364248 4196
rect 363104 4156 363110 4168
rect 364242 4156 364248 4168
rect 364300 4156 364306 4208
rect 368566 4156 368572 4208
rect 368624 4196 368630 4208
rect 369762 4196 369768 4208
rect 368624 4168 369768 4196
rect 368624 4156 368630 4168
rect 369762 4156 369768 4168
rect 369820 4156 369826 4208
rect 379606 4156 379612 4208
rect 379664 4196 379670 4208
rect 380802 4196 380808 4208
rect 379664 4168 380808 4196
rect 379664 4156 379670 4168
rect 380802 4156 380808 4168
rect 380860 4156 380866 4208
rect 401686 4156 401692 4208
rect 401744 4196 401750 4208
rect 402882 4196 402888 4208
rect 401744 4168 402888 4196
rect 401744 4156 401750 4168
rect 402882 4156 402888 4168
rect 402940 4156 402946 4208
rect 412726 4156 412732 4208
rect 412784 4196 412790 4208
rect 413922 4196 413928 4208
rect 412784 4168 413928 4196
rect 412784 4156 412790 4168
rect 413922 4156 413928 4168
rect 413980 4156 413986 4208
rect 59538 4088 59544 4140
rect 59596 4128 59602 4140
rect 253198 4128 253204 4140
rect 59596 4100 253204 4128
rect 59596 4088 59602 4100
rect 253198 4088 253204 4100
rect 253256 4088 253262 4140
rect 292942 4088 292948 4140
rect 293000 4128 293006 4140
rect 298002 4128 298008 4140
rect 293000 4100 298008 4128
rect 293000 4088 293006 4100
rect 298002 4088 298008 4100
rect 298060 4088 298066 4140
rect 316678 4088 316684 4140
rect 316736 4128 316742 4140
rect 440418 4128 440424 4140
rect 316736 4100 440424 4128
rect 316736 4088 316742 4100
rect 440418 4088 440424 4100
rect 440476 4088 440482 4140
rect 56226 4020 56232 4072
rect 56284 4060 56290 4072
rect 252646 4060 252652 4072
rect 56284 4032 252652 4060
rect 56284 4020 56290 4032
rect 252646 4020 252652 4032
rect 252704 4020 252710 4072
rect 317230 4020 317236 4072
rect 317288 4060 317294 4072
rect 443730 4060 443736 4072
rect 317288 4032 443736 4060
rect 317288 4020 317294 4032
rect 443730 4020 443736 4032
rect 443788 4020 443794 4072
rect 451366 4020 451372 4072
rect 451424 4060 451430 4072
rect 452562 4060 452568 4072
rect 451424 4032 452568 4060
rect 451424 4020 451430 4032
rect 452562 4020 452568 4032
rect 452620 4020 452626 4072
rect 52914 3952 52920 4004
rect 52972 3992 52978 4004
rect 252094 3992 252100 4004
rect 52972 3964 252100 3992
rect 52972 3952 52978 3964
rect 252094 3952 252100 3964
rect 252152 3952 252158 4004
rect 284754 3952 284760 4004
rect 284812 3992 284818 4004
rect 290734 3992 290740 4004
rect 284812 3964 290740 3992
rect 284812 3952 284818 3964
rect 290734 3952 290740 3964
rect 290792 3952 290798 4004
rect 317782 3952 317788 4004
rect 317840 3992 317846 4004
rect 447042 3992 447048 4004
rect 317840 3964 447048 3992
rect 317840 3952 317846 3964
rect 447042 3952 447048 3964
rect 447100 3952 447106 4004
rect 453666 3992 453672 4004
rect 451246 3964 453672 3992
rect 25314 3884 25320 3936
rect 25372 3924 25378 3936
rect 28258 3924 28264 3936
rect 25372 3896 28264 3924
rect 25372 3884 25378 3896
rect 28258 3884 28264 3896
rect 28316 3884 28322 3936
rect 49602 3884 49608 3936
rect 49660 3924 49666 3936
rect 251542 3924 251548 3936
rect 49660 3896 251548 3924
rect 49660 3884 49666 3896
rect 251542 3884 251548 3896
rect 251600 3884 251606 3936
rect 286962 3884 286968 3936
rect 287020 3924 287026 3936
rect 291378 3924 291384 3936
rect 287020 3896 291384 3924
rect 287020 3884 287026 3896
rect 291378 3884 291384 3896
rect 291436 3884 291442 3936
rect 292758 3884 292764 3936
rect 292816 3924 292822 3936
rect 296898 3924 296904 3936
rect 292816 3896 296904 3924
rect 292816 3884 292822 3896
rect 296898 3884 296904 3896
rect 296956 3884 296962 3936
rect 318334 3884 318340 3936
rect 318392 3924 318398 3936
rect 450354 3924 450360 3936
rect 318392 3896 450360 3924
rect 318392 3884 318398 3896
rect 450354 3884 450360 3896
rect 450412 3884 450418 3936
rect 46290 3816 46296 3868
rect 46348 3856 46354 3868
rect 250990 3856 250996 3868
rect 46348 3828 250996 3856
rect 46348 3816 46354 3828
rect 250990 3816 250996 3828
rect 251048 3816 251054 3868
rect 283650 3816 283656 3868
rect 283708 3856 283714 3868
rect 290550 3856 290556 3868
rect 283708 3828 290556 3856
rect 283708 3816 283714 3828
rect 290550 3816 290556 3828
rect 290608 3816 290614 3868
rect 318886 3816 318892 3868
rect 318944 3856 318950 3868
rect 451246 3856 451274 3964
rect 453666 3952 453672 3964
rect 453724 3952 453730 4004
rect 318944 3828 451274 3856
rect 318944 3816 318950 3828
rect 42978 3748 42984 3800
rect 43036 3788 43042 3800
rect 250438 3788 250444 3800
rect 43036 3760 250444 3788
rect 43036 3748 43042 3760
rect 250438 3748 250444 3760
rect 250496 3748 250502 3800
rect 281442 3748 281448 3800
rect 281500 3788 281506 3800
rect 290182 3788 290188 3800
rect 281500 3760 290188 3788
rect 281500 3748 281506 3760
rect 290182 3748 290188 3760
rect 290240 3748 290246 3800
rect 319438 3748 319444 3800
rect 319496 3788 319502 3800
rect 456978 3788 456984 3800
rect 319496 3760 456984 3788
rect 319496 3748 319502 3760
rect 456978 3748 456984 3760
rect 457036 3748 457042 3800
rect 41874 3680 41880 3732
rect 41932 3720 41938 3732
rect 250254 3720 250260 3732
rect 41932 3692 250260 3720
rect 41932 3680 41938 3692
rect 250254 3680 250260 3692
rect 250312 3680 250318 3732
rect 278130 3680 278136 3732
rect 278188 3720 278194 3732
rect 289630 3720 289636 3732
rect 278188 3692 289636 3720
rect 278188 3680 278194 3692
rect 289630 3680 289636 3692
rect 289688 3680 289694 3732
rect 319990 3680 319996 3732
rect 320048 3720 320054 3732
rect 460290 3720 460296 3732
rect 320048 3692 460296 3720
rect 320048 3680 320054 3692
rect 460290 3680 460296 3692
rect 460348 3680 460354 3732
rect 38562 3612 38568 3664
rect 38620 3652 38626 3664
rect 38620 3624 44220 3652
rect 38620 3612 38626 3624
rect 33042 3544 33048 3596
rect 33100 3584 33106 3596
rect 35158 3584 35164 3596
rect 33100 3556 35164 3584
rect 33100 3544 33106 3556
rect 35158 3544 35164 3556
rect 35216 3544 35222 3596
rect 42794 3544 42800 3596
rect 42852 3584 42858 3596
rect 44082 3584 44088 3596
rect 42852 3556 44088 3584
rect 42852 3544 42858 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44192 3584 44220 3624
rect 44266 3612 44272 3664
rect 44324 3652 44330 3664
rect 249518 3652 249524 3664
rect 44324 3624 249524 3652
rect 44324 3612 44330 3624
rect 249518 3612 249524 3624
rect 249576 3612 249582 3664
rect 274818 3612 274824 3664
rect 274876 3652 274882 3664
rect 288618 3652 288624 3664
rect 274876 3624 288624 3652
rect 274876 3612 274882 3624
rect 288618 3612 288624 3624
rect 288676 3612 288682 3664
rect 292390 3612 292396 3664
rect 292448 3652 292454 3664
rect 294690 3652 294696 3664
rect 292448 3624 294696 3652
rect 292448 3612 292454 3624
rect 294690 3612 294696 3624
rect 294748 3612 294754 3664
rect 320542 3612 320548 3664
rect 320600 3652 320606 3664
rect 463602 3652 463608 3664
rect 320600 3624 463608 3652
rect 320600 3612 320606 3624
rect 463602 3612 463608 3624
rect 463660 3612 463666 3664
rect 467926 3612 467932 3664
rect 467984 3652 467990 3664
rect 469122 3652 469128 3664
rect 467984 3624 469128 3652
rect 467984 3612 467990 3624
rect 469122 3612 469128 3624
rect 469180 3612 469186 3664
rect 478966 3612 478972 3664
rect 479024 3652 479030 3664
rect 480162 3652 480168 3664
rect 479024 3624 480168 3652
rect 479024 3612 479030 3624
rect 480162 3612 480168 3624
rect 480220 3612 480226 3664
rect 484486 3612 484492 3664
rect 484544 3652 484550 3664
rect 485682 3652 485688 3664
rect 484544 3624 485688 3652
rect 484544 3612 484550 3624
rect 485682 3612 485688 3624
rect 485740 3612 485746 3664
rect 495526 3612 495532 3664
rect 495584 3652 495590 3664
rect 496722 3652 496728 3664
rect 495584 3624 496728 3652
rect 495584 3612 495590 3624
rect 496722 3612 496728 3624
rect 496780 3612 496786 3664
rect 523126 3612 523132 3664
rect 523184 3652 523190 3664
rect 524322 3652 524328 3664
rect 523184 3624 524328 3652
rect 523184 3612 523190 3624
rect 524322 3612 524328 3624
rect 524380 3612 524386 3664
rect 528646 3612 528652 3664
rect 528704 3652 528710 3664
rect 529842 3652 529848 3664
rect 528704 3624 529848 3652
rect 528704 3612 528710 3624
rect 529842 3612 529848 3624
rect 529900 3612 529906 3664
rect 534166 3612 534172 3664
rect 534224 3652 534230 3664
rect 535362 3652 535368 3664
rect 534224 3624 535368 3652
rect 534224 3612 534230 3624
rect 535362 3612 535368 3624
rect 535420 3612 535426 3664
rect 552658 3612 552664 3664
rect 552716 3652 552722 3664
rect 555234 3652 555240 3664
rect 552716 3624 555240 3652
rect 552716 3612 552722 3624
rect 555234 3612 555240 3624
rect 555292 3612 555298 3664
rect 249978 3584 249984 3596
rect 44192 3556 249984 3584
rect 249978 3544 249984 3556
rect 250036 3544 250042 3596
rect 271506 3544 271512 3596
rect 271564 3584 271570 3596
rect 288894 3584 288900 3596
rect 271564 3556 288900 3584
rect 271564 3544 271570 3556
rect 288894 3544 288900 3556
rect 288952 3544 288958 3596
rect 292206 3544 292212 3596
rect 292264 3584 292270 3596
rect 293586 3584 293592 3596
rect 292264 3556 293592 3584
rect 292264 3544 292270 3556
rect 293586 3544 293592 3556
rect 293644 3544 293650 3596
rect 336918 3544 336924 3596
rect 336976 3584 336982 3596
rect 562962 3584 562968 3596
rect 336976 3556 562968 3584
rect 336976 3544 336982 3556
rect 562962 3544 562968 3556
rect 563020 3544 563026 3596
rect 34146 3476 34152 3528
rect 34204 3516 34210 3528
rect 248966 3516 248972 3528
rect 34204 3488 248972 3516
rect 34204 3476 34210 3488
rect 248966 3476 248972 3488
rect 249024 3476 249030 3528
rect 268194 3476 268200 3528
rect 268252 3516 268258 3528
rect 287974 3516 287980 3528
rect 268252 3488 287980 3516
rect 268252 3476 268258 3488
rect 287974 3476 287980 3488
rect 288032 3476 288038 3528
rect 288066 3476 288072 3528
rect 288124 3516 288130 3528
rect 291470 3516 291476 3528
rect 288124 3488 291476 3516
rect 288124 3476 288130 3488
rect 291470 3476 291476 3488
rect 291528 3476 291534 3528
rect 313274 3476 313280 3528
rect 313332 3516 313338 3528
rect 314562 3516 314568 3528
rect 313332 3488 314568 3516
rect 313332 3476 313338 3488
rect 314562 3476 314568 3488
rect 314620 3476 314626 3528
rect 321278 3476 321284 3528
rect 321336 3516 321342 3528
rect 466914 3516 466920 3528
rect 321336 3488 466920 3516
rect 321336 3476 321342 3488
rect 466914 3476 466920 3488
rect 466972 3476 466978 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 491202 3516 491208 3528
rect 489972 3488 491208 3516
rect 489972 3476 489978 3488
rect 491202 3476 491208 3488
rect 491260 3476 491266 3528
rect 500954 3476 500960 3528
rect 501012 3516 501018 3528
rect 502242 3516 502248 3528
rect 501012 3488 502248 3516
rect 501012 3476 501018 3488
rect 502242 3476 502248 3488
rect 502300 3476 502306 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507762 3516 507768 3528
rect 506532 3488 507768 3516
rect 506532 3476 506538 3488
rect 507762 3476 507768 3488
rect 507820 3476 507826 3528
rect 511994 3476 512000 3528
rect 512052 3516 512058 3528
rect 513282 3516 513288 3528
rect 512052 3488 513288 3516
rect 512052 3476 512058 3488
rect 513282 3476 513288 3488
rect 513340 3476 513346 3528
rect 517514 3476 517520 3528
rect 517572 3516 517578 3528
rect 518802 3516 518808 3528
rect 517572 3488 518808 3516
rect 517572 3476 517578 3488
rect 518802 3476 518808 3488
rect 518860 3476 518866 3528
rect 549898 3476 549904 3528
rect 549956 3516 549962 3528
rect 550818 3516 550824 3528
rect 549956 3488 550824 3516
rect 549956 3476 549962 3488
rect 550818 3476 550824 3488
rect 550876 3476 550882 3528
rect 29730 3408 29736 3460
rect 29788 3448 29794 3460
rect 241422 3448 241428 3460
rect 29788 3420 241428 3448
rect 29788 3408 29794 3420
rect 241422 3408 241428 3420
rect 241480 3408 241486 3460
rect 241514 3408 241520 3460
rect 241572 3448 241578 3460
rect 242802 3448 242808 3460
rect 241572 3420 242808 3448
rect 241572 3408 241578 3420
rect 242802 3408 242808 3420
rect 242860 3408 242866 3460
rect 264882 3408 264888 3460
rect 264940 3448 264946 3460
rect 287514 3448 287520 3460
rect 264940 3420 287520 3448
rect 264940 3408 264946 3420
rect 287514 3408 287520 3420
rect 287572 3408 287578 3460
rect 290274 3408 290280 3460
rect 290332 3448 290338 3460
rect 291746 3448 291752 3460
rect 290332 3420 291752 3448
rect 290332 3408 290338 3420
rect 291746 3408 291752 3420
rect 291804 3408 291810 3460
rect 293494 3408 293500 3460
rect 293552 3448 293558 3460
rect 301314 3448 301320 3460
rect 293552 3420 301320 3448
rect 293552 3408 293558 3420
rect 301314 3408 301320 3420
rect 301372 3408 301378 3460
rect 340874 3408 340880 3460
rect 340932 3448 340938 3460
rect 342162 3448 342168 3460
rect 340932 3420 342168 3448
rect 340932 3408 340938 3420
rect 342162 3408 342168 3420
rect 342220 3408 342226 3460
rect 342254 3408 342260 3460
rect 342312 3448 342318 3460
rect 561858 3448 561864 3460
rect 342312 3420 561864 3448
rect 342312 3408 342318 3420
rect 561858 3408 561864 3420
rect 561916 3408 561922 3460
rect 37458 3340 37464 3392
rect 37516 3380 37522 3392
rect 44266 3380 44272 3392
rect 37516 3352 44272 3380
rect 37516 3340 37522 3352
rect 44266 3340 44272 3352
rect 44324 3340 44330 3392
rect 53834 3340 53840 3392
rect 53892 3380 53898 3392
rect 55122 3380 55128 3392
rect 53892 3352 55128 3380
rect 53892 3340 53898 3352
rect 55122 3340 55128 3352
rect 55180 3340 55186 3392
rect 59354 3340 59360 3392
rect 59412 3380 59418 3392
rect 60642 3380 60648 3392
rect 59412 3352 60648 3380
rect 59412 3340 59418 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 62850 3340 62856 3392
rect 62908 3380 62914 3392
rect 253750 3380 253756 3392
rect 62908 3352 253756 3380
rect 62908 3340 62914 3352
rect 253750 3340 253756 3352
rect 253808 3340 253814 3392
rect 292574 3340 292580 3392
rect 292632 3380 292638 3392
rect 295794 3380 295800 3392
rect 292632 3352 295800 3380
rect 292632 3340 292638 3352
rect 295794 3340 295800 3352
rect 295852 3340 295858 3392
rect 316126 3340 316132 3392
rect 316184 3380 316190 3392
rect 316184 3352 434668 3380
rect 316184 3340 316190 3352
rect 75914 3272 75920 3324
rect 75972 3312 75978 3324
rect 77202 3312 77208 3324
rect 75972 3284 77208 3312
rect 75972 3272 75978 3284
rect 77202 3272 77208 3284
rect 77260 3272 77266 3324
rect 81434 3272 81440 3324
rect 81492 3312 81498 3324
rect 82722 3312 82728 3324
rect 81492 3284 82728 3312
rect 81492 3272 81498 3284
rect 82722 3272 82728 3284
rect 82780 3272 82786 3324
rect 92474 3272 92480 3324
rect 92532 3312 92538 3324
rect 93762 3312 93768 3324
rect 92532 3284 93768 3312
rect 92532 3272 92538 3284
rect 93762 3272 93768 3284
rect 93820 3272 93826 3324
rect 97994 3272 98000 3324
rect 98052 3312 98058 3324
rect 99282 3312 99288 3324
rect 98052 3284 99288 3312
rect 98052 3272 98058 3284
rect 99282 3272 99288 3284
rect 99340 3272 99346 3324
rect 103514 3272 103520 3324
rect 103572 3312 103578 3324
rect 104802 3312 104808 3324
rect 103572 3284 104808 3312
rect 103572 3272 103578 3284
rect 104802 3272 104808 3284
rect 104860 3272 104866 3324
rect 109034 3272 109040 3324
rect 109092 3312 109098 3324
rect 110322 3312 110328 3324
rect 109092 3284 110328 3312
rect 109092 3272 109098 3284
rect 110322 3272 110328 3284
rect 110380 3272 110386 3324
rect 125594 3272 125600 3324
rect 125652 3312 125658 3324
rect 126882 3312 126888 3324
rect 125652 3284 126888 3312
rect 125652 3272 125658 3284
rect 126882 3272 126888 3284
rect 126940 3272 126946 3324
rect 132402 3272 132408 3324
rect 132460 3312 132466 3324
rect 265526 3312 265532 3324
rect 132460 3284 265532 3312
rect 132460 3272 132466 3284
rect 265526 3272 265532 3284
rect 265584 3272 265590 3324
rect 315574 3272 315580 3324
rect 315632 3312 315638 3324
rect 433794 3312 433800 3324
rect 315632 3284 433800 3312
rect 315632 3272 315638 3284
rect 433794 3272 433800 3284
rect 433852 3272 433858 3324
rect 434640 3312 434668 3352
rect 434714 3340 434720 3392
rect 434772 3380 434778 3392
rect 436002 3380 436008 3392
rect 434772 3352 436008 3380
rect 434772 3340 434778 3352
rect 436002 3340 436008 3352
rect 436060 3340 436066 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 456886 3340 456892 3392
rect 456944 3380 456950 3392
rect 458082 3380 458088 3392
rect 456944 3352 458088 3380
rect 456944 3340 456950 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 550726 3340 550732 3392
rect 550784 3380 550790 3392
rect 551922 3380 551928 3392
rect 550784 3352 551928 3380
rect 550784 3340 550790 3352
rect 551922 3340 551928 3352
rect 551980 3340 551986 3392
rect 437106 3312 437112 3324
rect 434640 3284 437112 3312
rect 437106 3272 437112 3284
rect 437164 3272 437170 3324
rect 135714 3204 135720 3256
rect 135772 3244 135778 3256
rect 265894 3244 265900 3256
rect 135772 3216 265900 3244
rect 135772 3204 135778 3216
rect 265894 3204 265900 3216
rect 265952 3204 265958 3256
rect 315022 3204 315028 3256
rect 315080 3244 315086 3256
rect 315080 3216 412634 3244
rect 315080 3204 315086 3216
rect 142154 3136 142160 3188
rect 142212 3176 142218 3188
rect 143442 3176 143448 3188
rect 142212 3148 143448 3176
rect 142212 3136 142218 3148
rect 143442 3136 143448 3148
rect 143500 3136 143506 3188
rect 158714 3136 158720 3188
rect 158772 3176 158778 3188
rect 160002 3176 160008 3188
rect 158772 3148 160008 3176
rect 158772 3136 158778 3148
rect 160002 3136 160008 3148
rect 160060 3136 160066 3188
rect 175274 3136 175280 3188
rect 175332 3176 175338 3188
rect 176562 3176 176568 3188
rect 175332 3148 176568 3176
rect 175332 3136 175338 3148
rect 176562 3136 176568 3148
rect 176620 3136 176626 3188
rect 186314 3136 186320 3188
rect 186372 3176 186378 3188
rect 187602 3176 187608 3188
rect 186372 3148 187608 3176
rect 186372 3136 186378 3148
rect 187602 3136 187608 3148
rect 187660 3136 187666 3188
rect 191834 3136 191840 3188
rect 191892 3176 191898 3188
rect 193122 3176 193128 3188
rect 191892 3148 193128 3176
rect 191892 3136 191898 3148
rect 193122 3136 193128 3148
rect 193180 3136 193186 3188
rect 208394 3136 208400 3188
rect 208452 3176 208458 3188
rect 209682 3176 209688 3188
rect 208452 3148 209688 3176
rect 208452 3136 208458 3148
rect 209682 3136 209688 3148
rect 209740 3136 209746 3188
rect 219434 3136 219440 3188
rect 219492 3176 219498 3188
rect 220722 3176 220728 3188
rect 219492 3148 220728 3176
rect 219492 3136 219498 3148
rect 220722 3136 220728 3148
rect 220780 3136 220786 3188
rect 224954 3136 224960 3188
rect 225012 3176 225018 3188
rect 226242 3176 226248 3188
rect 225012 3148 226248 3176
rect 225012 3136 225018 3148
rect 226242 3136 226248 3148
rect 226300 3136 226306 3188
rect 241422 3136 241428 3188
rect 241480 3176 241486 3188
rect 248230 3176 248236 3188
rect 241480 3148 248236 3176
rect 241480 3136 241486 3148
rect 248230 3136 248236 3148
rect 248288 3136 248294 3188
rect 289170 3136 289176 3188
rect 289228 3176 289234 3188
rect 291562 3176 291568 3188
rect 289228 3148 291568 3176
rect 289228 3136 289234 3148
rect 291562 3136 291568 3148
rect 291620 3136 291626 3188
rect 336734 3136 336740 3188
rect 336792 3176 336798 3188
rect 342254 3176 342260 3188
rect 336792 3148 342260 3176
rect 336792 3136 336798 3148
rect 342254 3136 342260 3148
rect 342312 3136 342318 3188
rect 357434 3136 357440 3188
rect 357492 3176 357498 3188
rect 358722 3176 358728 3188
rect 357492 3148 358728 3176
rect 357492 3136 357498 3148
rect 358722 3136 358728 3148
rect 358780 3136 358786 3188
rect 373994 3136 374000 3188
rect 374052 3176 374058 3188
rect 375282 3176 375288 3188
rect 374052 3148 375288 3176
rect 374052 3136 374058 3148
rect 375282 3136 375288 3148
rect 375340 3136 375346 3188
rect 385034 3136 385040 3188
rect 385092 3176 385098 3188
rect 386322 3176 386328 3188
rect 385092 3148 386328 3176
rect 385092 3136 385098 3148
rect 386322 3136 386328 3148
rect 386380 3136 386386 3188
rect 390554 3136 390560 3188
rect 390612 3176 390618 3188
rect 391842 3176 391848 3188
rect 390612 3148 391848 3176
rect 390612 3136 390618 3148
rect 391842 3136 391848 3148
rect 391900 3136 391906 3188
rect 396074 3136 396080 3188
rect 396132 3176 396138 3188
rect 397362 3176 397368 3188
rect 396132 3148 397368 3176
rect 396132 3136 396138 3148
rect 397362 3136 397368 3148
rect 397420 3136 397426 3188
rect 407114 3136 407120 3188
rect 407172 3176 407178 3188
rect 408402 3176 408408 3188
rect 407172 3148 408408 3176
rect 407172 3136 407178 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 412606 3176 412634 3216
rect 418154 3204 418160 3256
rect 418212 3244 418218 3256
rect 419442 3244 419448 3256
rect 418212 3216 419448 3244
rect 418212 3204 418218 3216
rect 419442 3204 419448 3216
rect 419500 3204 419506 3256
rect 423674 3204 423680 3256
rect 423732 3244 423738 3256
rect 424962 3244 424968 3256
rect 423732 3216 424968 3244
rect 423732 3204 423738 3216
rect 424962 3204 424968 3216
rect 425020 3204 425026 3256
rect 430482 3176 430488 3188
rect 412606 3148 430488 3176
rect 430482 3136 430488 3148
rect 430540 3136 430546 3188
rect 27522 3000 27528 3052
rect 27580 3040 27586 3052
rect 32398 3040 32404 3052
rect 27580 3012 32404 3040
rect 27580 3000 27586 3012
rect 32398 3000 32404 3012
rect 32456 3000 32462 3052
rect 136634 2728 136640 2780
rect 136692 2768 136698 2780
rect 137922 2768 137928 2780
rect 136692 2740 137928 2768
rect 136692 2728 136698 2740
rect 137922 2728 137928 2740
rect 137980 2728 137986 2780
rect 335354 2592 335360 2644
rect 335412 2632 335418 2644
rect 336642 2632 336648 2644
rect 335412 2604 336648 2632
rect 335412 2592 335418 2604
rect 336642 2592 336648 2604
rect 336700 2592 336706 2644
rect 329834 2388 329840 2440
rect 329892 2428 329898 2440
rect 331122 2428 331128 2440
rect 329892 2400 331128 2428
rect 329892 2388 329898 2400
rect 331122 2388 331128 2400
rect 331180 2388 331186 2440
rect 20714 2320 20720 2372
rect 20772 2360 20778 2372
rect 22002 2360 22008 2372
rect 20772 2332 22008 2360
rect 20772 2320 20778 2332
rect 22002 2320 22008 2332
rect 22060 2320 22066 2372
rect 539594 1232 539600 1284
rect 539652 1272 539658 1284
rect 540882 1272 540888 1284
rect 539652 1244 540888 1272
rect 539652 1232 539658 1244
rect 540882 1232 540888 1244
rect 540940 1232 540946 1284
rect 545114 1232 545120 1284
rect 545172 1272 545178 1284
rect 546402 1272 546408 1284
rect 545172 1244 546408 1272
rect 545172 1232 545178 1244
rect 546402 1232 546408 1244
rect 546460 1232 546466 1284
rect 556154 1232 556160 1284
rect 556212 1272 556218 1284
rect 557442 1272 557448 1284
rect 556212 1244 557448 1272
rect 556212 1232 556218 1244
rect 557442 1232 557448 1244
rect 557500 1232 557506 1284
<< via1 >>
rect 88340 702992 88392 703044
rect 89536 702992 89588 703044
rect 309140 700884 309192 700936
rect 364800 700884 364852 700936
rect 313280 700816 313332 700868
rect 397184 700816 397236 700868
rect 317420 700748 317472 700800
rect 413376 700748 413428 700800
rect 321560 700680 321612 700732
rect 429568 700680 429620 700732
rect 327080 700612 327132 700664
rect 461952 700612 462004 700664
rect 331312 700544 331364 700596
rect 478144 700544 478196 700596
rect 295340 700476 295392 700528
rect 300032 700476 300084 700528
rect 335360 700476 335412 700528
rect 494336 700476 494388 700528
rect 339500 700408 339552 700460
rect 526720 700408 526772 700460
rect 299480 700340 299532 700392
rect 332416 700340 332468 700392
rect 343640 700340 343692 700392
rect 542912 700340 542964 700392
rect 267648 700272 267700 700324
rect 279424 700272 279476 700324
rect 305000 700272 305052 700324
rect 348608 700272 348660 700324
rect 349160 700272 349212 700324
rect 559104 700272 559156 700324
rect 23480 697552 23532 697604
rect 24768 697552 24820 697604
rect 2780 680552 2832 680604
rect 4804 680552 4856 680604
rect 353944 680348 353996 680400
rect 580172 680348 580224 680400
rect 360844 667904 360896 667956
rect 580172 667904 580224 667956
rect 367744 641724 367796 641776
rect 579896 641724 579948 641776
rect 3608 629280 3660 629332
rect 35164 629280 35216 629332
rect 377404 627920 377456 627972
rect 579896 627920 579948 627972
rect 3332 615476 3384 615528
rect 22744 615476 22796 615528
rect 509884 615476 509936 615528
rect 580172 615476 580224 615528
rect 3332 603100 3384 603152
rect 14464 603100 14516 603152
rect 3332 576852 3384 576904
rect 7564 576852 7616 576904
rect 359464 561688 359516 561740
rect 580172 561688 580224 561740
rect 364984 535440 365036 535492
rect 580172 535440 580224 535492
rect 3332 525784 3384 525836
rect 61384 525784 61436 525836
rect 374644 522996 374696 523048
rect 580172 522996 580224 523048
rect 3332 513340 3384 513392
rect 25504 513340 25556 513392
rect 356704 509260 356756 509312
rect 579620 509260 579672 509312
rect 2964 499536 3016 499588
rect 17224 499536 17276 499588
rect 3240 474036 3292 474088
rect 8944 474036 8996 474088
rect 355324 456764 355376 456816
rect 580172 456764 580224 456816
rect 373264 430584 373316 430636
rect 579804 430584 579856 430636
rect 2964 422288 3016 422340
rect 180064 422288 180116 422340
rect 381544 416780 381596 416832
rect 579620 416780 579672 416832
rect 3332 409844 3384 409896
rect 26884 409844 26936 409896
rect 363604 404336 363656 404388
rect 580172 404336 580224 404388
rect 2964 396040 3016 396092
rect 18604 396040 18656 396092
rect 3332 371220 3384 371272
rect 10324 371220 10376 371272
rect 354036 364352 354088 364404
rect 580172 364352 580224 364404
rect 371884 324300 371936 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 224224 318792 224276 318844
rect 378784 311856 378836 311908
rect 580172 311856 580224 311908
rect 3332 306348 3384 306400
rect 28264 306348 28316 306400
rect 3332 292544 3384 292596
rect 21364 292544 21416 292596
rect 369124 271872 369176 271924
rect 579988 271872 580040 271924
rect 3332 267724 3384 267776
rect 13084 267724 13136 267776
rect 218060 263508 218112 263560
rect 278688 263508 278740 263560
rect 202880 263440 202932 263492
rect 274272 263440 274324 263492
rect 169760 263372 169812 263424
rect 269856 263372 269908 263424
rect 153200 263304 153252 263356
rect 265440 263304 265492 263356
rect 138020 263236 138072 263288
rect 261024 263236 261076 263288
rect 104900 263168 104952 263220
rect 256608 263168 256660 263220
rect 88340 263100 88392 263152
rect 252192 263100 252244 263152
rect 73160 263032 73212 263084
rect 247776 263032 247828 263084
rect 40040 262964 40092 263016
rect 243360 262964 243412 263016
rect 282920 262964 282972 263016
rect 291936 262964 291988 263016
rect 23480 262896 23532 262948
rect 238944 262896 238996 262948
rect 279424 262896 279476 262948
rect 287520 262896 287572 262948
rect 8300 262828 8352 262880
rect 234528 262828 234580 262880
rect 234620 262828 234672 262880
rect 283104 262828 283156 262880
rect 354128 259428 354180 259480
rect 580172 259428 580224 259480
rect 4804 258000 4856 258052
rect 230388 258000 230440 258052
rect 353300 258000 353352 258052
rect 580172 258000 580224 258052
rect 3424 255212 3476 255264
rect 230388 255212 230440 255264
rect 3516 251132 3568 251184
rect 230388 251132 230440 251184
rect 353300 251132 353352 251184
rect 360844 251132 360896 251184
rect 353300 248344 353352 248396
rect 367744 248344 367796 248396
rect 35164 246984 35216 247036
rect 229652 246984 229704 247036
rect 353300 244196 353352 244248
rect 377404 244196 377456 244248
rect 22744 242836 22796 242888
rect 229284 242836 229336 242888
rect 14464 240048 14516 240100
rect 230020 240048 230072 240100
rect 353300 240048 353352 240100
rect 509884 240048 509936 240100
rect 353300 237328 353352 237380
rect 580356 237328 580408 237380
rect 7564 235900 7616 235952
rect 230204 235900 230256 235952
rect 353300 233180 353352 233232
rect 580448 233180 580500 233232
rect 3608 231752 3660 231804
rect 230388 231752 230440 231804
rect 353300 230392 353352 230444
rect 359464 230392 359516 230444
rect 3700 227672 3752 227724
rect 230388 227672 230440 227724
rect 353300 226244 353352 226296
rect 364984 226244 365036 226296
rect 61384 224884 61436 224936
rect 229652 224884 229704 224936
rect 353300 223524 353352 223576
rect 374644 223524 374696 223576
rect 25504 220736 25556 220788
rect 230388 220736 230440 220788
rect 353944 219444 353996 219496
rect 580172 219444 580224 219496
rect 353300 219376 353352 219428
rect 356704 219376 356756 219428
rect 17224 216588 17276 216640
rect 230388 216588 230440 216640
rect 353300 215228 353352 215280
rect 580540 215228 580592 215280
rect 8944 212440 8996 212492
rect 230388 212440 230440 212492
rect 353300 212440 353352 212492
rect 580632 212440 580684 212492
rect 3792 209720 3844 209772
rect 229652 209720 229704 209772
rect 353300 208156 353352 208208
rect 355324 208156 355376 208208
rect 3884 205572 3936 205624
rect 229468 205572 229520 205624
rect 353300 205572 353352 205624
rect 373264 205572 373316 205624
rect 180064 201424 180116 201476
rect 230388 201424 230440 201476
rect 353300 201424 353352 201476
rect 381544 201424 381596 201476
rect 353300 198636 353352 198688
rect 363604 198636 363656 198688
rect 26884 197276 26936 197328
rect 229836 197276 229888 197328
rect 353300 194488 353352 194540
rect 580724 194488 580776 194540
rect 18604 193128 18656 193180
rect 230388 193128 230440 193180
rect 10324 190408 10376 190460
rect 230388 190408 230440 190460
rect 353300 187620 353352 187672
rect 580816 187620 580868 187672
rect 3976 186260 4028 186312
rect 230388 186260 230440 186312
rect 353300 183472 353352 183524
rect 371884 183472 371936 183524
rect 4068 182112 4120 182164
rect 229836 182112 229888 182164
rect 353300 180752 353352 180804
rect 378784 180752 378836 180804
rect 354036 179392 354088 179444
rect 579620 179392 579672 179444
rect 224224 177964 224276 178016
rect 230388 177964 230440 178016
rect 353300 176604 353352 176656
rect 580908 176604 580960 176656
rect 28264 175176 28316 175228
rect 230388 175176 230440 175228
rect 353300 173816 353352 173868
rect 369124 173816 369176 173868
rect 21364 171028 21416 171080
rect 230388 171028 230440 171080
rect 13084 166948 13136 167000
rect 230388 166948 230440 167000
rect 353300 166948 353352 167000
rect 580264 166948 580316 167000
rect 3332 162800 3384 162852
rect 230388 162800 230440 162852
rect 353300 162800 353352 162852
rect 580356 162800 580408 162852
rect 3424 160012 3476 160064
rect 230388 160012 230440 160064
rect 3516 155864 3568 155916
rect 229284 155864 229336 155916
rect 353300 155864 353352 155916
rect 580448 155864 580500 155916
rect 353944 153212 353996 153264
rect 579620 153212 579672 153264
rect 3608 151716 3660 151768
rect 230388 151716 230440 151768
rect 353300 151716 353352 151768
rect 580540 151716 580592 151768
rect 3700 147568 3752 147620
rect 230388 147568 230440 147620
rect 3792 144848 3844 144900
rect 230020 144848 230072 144900
rect 353300 144848 353352 144900
rect 580632 144848 580684 144900
rect 353300 140768 353352 140820
rect 580172 140768 580224 140820
rect 3424 140700 3476 140752
rect 230388 140700 230440 140752
rect 3424 136552 3476 136604
rect 229652 136552 229704 136604
rect 3608 128324 3660 128376
rect 230388 128324 230440 128376
rect 354220 128256 354272 128308
rect 580172 128256 580224 128308
rect 3516 115948 3568 116000
rect 230388 115948 230440 116000
rect 353944 114452 353996 114504
rect 580172 114452 580224 114504
rect 3148 113092 3200 113144
rect 229744 113092 229796 113144
rect 3424 104864 3476 104916
rect 230388 104864 230440 104916
rect 354588 102076 354640 102128
rect 579988 102076 580040 102128
rect 247684 97928 247736 97980
rect 248512 97928 248564 97980
rect 286324 97928 286376 97980
rect 287336 97928 287388 97980
rect 303896 97928 303948 97980
rect 307116 97928 307168 97980
rect 246948 97860 247000 97912
rect 249984 97860 250036 97912
rect 276756 97860 276808 97912
rect 277768 97860 277820 97912
rect 284944 97860 284996 97912
rect 287152 97860 287204 97912
rect 332968 97860 333020 97912
rect 338764 97860 338816 97912
rect 244924 97792 244976 97844
rect 255688 97792 255740 97844
rect 282276 97792 282328 97844
rect 288808 97792 288860 97844
rect 294144 97792 294196 97844
rect 300308 97792 300360 97844
rect 334624 97792 334676 97844
rect 337476 97792 337528 97844
rect 235264 97724 235316 97776
rect 249248 97724 249300 97776
rect 294880 97724 294932 97776
rect 301780 97724 301832 97776
rect 325792 97724 325844 97776
rect 339040 97724 339092 97776
rect 243544 97656 243596 97708
rect 266176 97656 266228 97708
rect 293960 97656 294012 97708
rect 300860 97656 300912 97708
rect 316408 97656 316460 97708
rect 326344 97656 326396 97708
rect 330760 97656 330812 97708
rect 347044 97656 347096 97708
rect 242164 97588 242216 97640
rect 272248 97588 272300 97640
rect 278412 97588 278464 97640
rect 281080 97588 281132 97640
rect 295616 97588 295668 97640
rect 304540 97588 304592 97640
rect 321928 97588 321980 97640
rect 338856 97588 338908 97640
rect 239404 97520 239456 97572
rect 274456 97520 274508 97572
rect 279884 97520 279936 97572
rect 289360 97520 289412 97572
rect 294328 97520 294380 97572
rect 303620 97520 303672 97572
rect 322480 97520 322532 97572
rect 341524 97520 341576 97572
rect 128360 97452 128412 97504
rect 264888 97452 264940 97504
rect 275284 97452 275336 97504
rect 285680 97452 285732 97504
rect 299296 97452 299348 97504
rect 322940 97452 322992 97504
rect 324688 97452 324740 97504
rect 342904 97452 342956 97504
rect 238024 97384 238076 97436
rect 281632 97384 281684 97436
rect 121460 97316 121512 97368
rect 263784 97316 263836 97368
rect 278044 97316 278096 97368
rect 288440 97384 288492 97436
rect 298192 97384 298244 97436
rect 324044 97384 324096 97436
rect 326896 97384 326948 97436
rect 345664 97384 345716 97436
rect 297088 97316 297140 97368
rect 320916 97316 320968 97368
rect 321376 97316 321428 97368
rect 349804 97316 349856 97368
rect 28264 97248 28316 97300
rect 247592 97248 247644 97300
rect 273996 97248 274048 97300
rect 264980 97180 265032 97232
rect 272800 97180 272852 97232
rect 278228 97248 278280 97300
rect 279056 97248 279108 97300
rect 286048 97248 286100 97300
rect 297640 97248 297692 97300
rect 323492 97248 323544 97300
rect 326436 97248 326488 97300
rect 475384 97248 475436 97300
rect 281540 97180 281592 97232
rect 283288 97180 283340 97232
rect 330208 97180 330260 97232
rect 338948 97180 339000 97232
rect 255964 97112 256016 97164
rect 258448 97112 258500 97164
rect 257436 96976 257488 97028
rect 259000 96976 259052 97028
rect 261024 96976 261076 97028
rect 261484 96976 261536 97028
rect 274180 96976 274232 97028
rect 277216 96976 277268 97028
rect 265164 96908 265216 96960
rect 265624 96908 265676 96960
rect 273628 96908 273680 96960
rect 274088 96908 274140 96960
rect 275100 96908 275152 96960
rect 275376 96908 275428 96960
rect 279608 96908 279660 96960
rect 280528 96908 280580 96960
rect 287152 96908 287204 96960
rect 287704 96908 287756 96960
rect 289176 96908 289228 96960
rect 289912 96908 289964 96960
rect 335728 96908 335780 96960
rect 337384 96908 337436 96960
rect 243636 96840 243688 96892
rect 247040 96840 247092 96892
rect 264244 96840 264296 96892
rect 266728 96840 266780 96892
rect 272524 96840 272576 96892
rect 274824 96840 274876 96892
rect 279700 96840 279752 96892
rect 286600 96840 286652 96892
rect 335360 96840 335412 96892
rect 340144 96840 340196 96892
rect 246396 96772 246448 96824
rect 247776 96772 247828 96824
rect 252928 96772 252980 96824
rect 253112 96772 253164 96824
rect 260932 96772 260984 96824
rect 261392 96772 261444 96824
rect 263692 96772 263744 96824
rect 264152 96772 264204 96824
rect 271144 96772 271196 96824
rect 271880 96772 271932 96824
rect 282184 96772 282236 96824
rect 284852 96772 284904 96824
rect 288624 96772 288676 96824
rect 289084 96772 289136 96824
rect 301136 96772 301188 96824
rect 302976 96772 303028 96824
rect 303620 96772 303672 96824
rect 304264 96772 304316 96824
rect 308128 96772 308180 96824
rect 309784 96772 309836 96824
rect 311992 96772 312044 96824
rect 315304 96772 315356 96824
rect 316960 96772 317012 96824
rect 318064 96772 318116 96824
rect 322940 96772 322992 96824
rect 323768 96772 323820 96824
rect 260104 96704 260156 96756
rect 262312 96704 262364 96756
rect 265624 96704 265676 96756
rect 267280 96704 267332 96756
rect 274088 96704 274140 96756
rect 275008 96704 275060 96756
rect 276664 96704 276716 96756
rect 277584 96704 277636 96756
rect 285864 96704 285916 96756
rect 287704 96704 287756 96756
rect 290464 96704 290516 96756
rect 300860 96704 300912 96756
rect 301504 96704 301556 96756
rect 318800 96704 318852 96756
rect 325056 96704 325108 96756
rect 246304 96636 246356 96688
rect 246948 96636 247000 96688
rect 257344 96636 257396 96688
rect 258080 96636 258132 96688
rect 269396 96568 269448 96620
rect 276112 96636 276164 96688
rect 279424 96636 279476 96688
rect 279884 96636 279936 96688
rect 283104 96636 283156 96688
rect 283472 96636 283524 96688
rect 283564 96636 283616 96688
rect 283656 96636 283708 96688
rect 284576 96636 284628 96688
rect 289084 96636 289136 96688
rect 290096 96636 290148 96688
rect 224960 96228 225012 96280
rect 278412 96228 278464 96280
rect 299848 96228 299900 96280
rect 338120 96228 338172 96280
rect 216680 96160 216732 96212
rect 279516 96160 279568 96212
rect 302608 96160 302660 96212
rect 354680 96160 354732 96212
rect 195980 96092 196032 96144
rect 269396 96092 269448 96144
rect 269488 96092 269540 96144
rect 269672 96092 269724 96144
rect 308680 96092 308732 96144
rect 390560 96092 390612 96144
rect 169760 96024 169812 96076
rect 271696 96024 271748 96076
rect 316040 96024 316092 96076
rect 434720 96024 434772 96076
rect 81440 95956 81492 96008
rect 257160 95956 257212 96008
rect 323032 95956 323084 96008
rect 477500 95956 477552 96008
rect 75920 95888 75972 95940
rect 256240 95888 256292 95940
rect 327448 95888 327500 95940
rect 503720 95888 503772 95940
rect 277860 95684 277912 95736
rect 278136 95684 278188 95736
rect 279424 95548 279476 95600
rect 279700 95548 279752 95600
rect 273996 95412 274048 95464
rect 274180 95412 274232 95464
rect 269120 95208 269172 95260
rect 269304 95208 269356 95260
rect 281632 95140 281684 95192
rect 282368 95140 282420 95192
rect 238760 94800 238812 94852
rect 281540 94800 281592 94852
rect 213920 94732 213972 94784
rect 278228 94732 278280 94784
rect 303160 94732 303212 94784
rect 357440 94732 357492 94784
rect 198740 94664 198792 94716
rect 276572 94664 276624 94716
rect 310704 94664 310756 94716
rect 402980 94664 403032 94716
rect 175280 94596 175332 94648
rect 264980 94596 265032 94648
rect 313648 94596 313700 94648
rect 420920 94596 420972 94648
rect 66260 94528 66312 94580
rect 254584 94528 254636 94580
rect 323584 94528 323636 94580
rect 480260 94528 480312 94580
rect 40040 94460 40092 94512
rect 250168 94460 250220 94512
rect 298744 94460 298796 94512
rect 331220 94460 331272 94512
rect 331312 94460 331364 94512
rect 527180 94460 527232 94512
rect 255320 94392 255372 94444
rect 255504 94392 255556 94444
rect 241520 93440 241572 93492
rect 283840 93440 283892 93492
rect 219440 93372 219492 93424
rect 280160 93372 280212 93424
rect 302976 93372 303028 93424
rect 346400 93372 346452 93424
rect 205640 93304 205692 93356
rect 276756 93304 276808 93356
rect 300952 93304 301004 93356
rect 345020 93304 345072 93356
rect 179420 93236 179472 93288
rect 273352 93236 273404 93288
rect 309784 93236 309836 93288
rect 387800 93236 387852 93288
rect 63500 93168 63552 93220
rect 254032 93168 254084 93220
rect 324136 93168 324188 93220
rect 484400 93168 484452 93220
rect 56600 93100 56652 93152
rect 253112 93100 253164 93152
rect 334072 93100 334124 93152
rect 543740 93100 543792 93152
rect 233240 92012 233292 92064
rect 281632 92012 281684 92064
rect 303712 92012 303764 92064
rect 361580 92012 361632 92064
rect 212540 91944 212592 91996
rect 278872 91944 278924 91996
rect 307944 91944 307996 91996
rect 386420 91944 386472 91996
rect 182180 91876 182232 91928
rect 273812 91876 273864 91928
rect 300400 91876 300452 91928
rect 340880 91876 340932 91928
rect 349804 91876 349856 91928
rect 467840 91876 467892 91928
rect 155960 91808 156012 91860
rect 269672 91808 269724 91860
rect 319168 91808 319220 91860
rect 454040 91808 454092 91860
rect 106280 91740 106332 91792
rect 261208 91740 261260 91792
rect 333520 91740 333572 91792
rect 539600 91740 539652 91792
rect 237380 90584 237432 90636
rect 283472 90584 283524 90636
rect 300032 90584 300084 90636
rect 339500 90584 339552 90636
rect 219532 90516 219584 90568
rect 279976 90516 280028 90568
rect 307024 90516 307076 90568
rect 362960 90516 363012 90568
rect 189080 90448 189132 90500
rect 274088 90448 274140 90500
rect 304172 90448 304224 90500
rect 364340 90448 364392 90500
rect 173900 90380 173952 90432
rect 272432 90380 272484 90432
rect 325240 90380 325292 90432
rect 489920 90380 489972 90432
rect 92480 90312 92532 90364
rect 257436 90312 257488 90364
rect 336280 90312 336332 90364
rect 556160 90312 556212 90364
rect 231860 89224 231912 89276
rect 282092 89224 282144 89276
rect 301412 89224 301464 89276
rect 347780 89224 347832 89276
rect 191840 89156 191892 89208
rect 275560 89156 275612 89208
rect 305368 89156 305420 89208
rect 371240 89156 371292 89208
rect 136640 89088 136692 89140
rect 266360 89088 266412 89140
rect 315304 89088 315356 89140
rect 411260 89088 411312 89140
rect 98000 89020 98052 89072
rect 259920 89020 259972 89072
rect 339040 89020 339092 89072
rect 494060 89020 494112 89072
rect 80060 88952 80112 89004
rect 256792 88952 256844 89004
rect 329840 88952 329892 89004
rect 517520 88952 517572 89004
rect 3332 88272 3384 88324
rect 230112 88272 230164 88324
rect 354496 88272 354548 88324
rect 580172 88272 580224 88324
rect 245844 87864 245896 87916
rect 284392 87864 284444 87916
rect 223580 87796 223632 87848
rect 280712 87796 280764 87848
rect 302056 87796 302108 87848
rect 351920 87796 351972 87848
rect 208400 87728 208452 87780
rect 278320 87728 278372 87780
rect 305920 87728 305972 87780
rect 374000 87728 374052 87780
rect 187700 87660 187752 87712
rect 272524 87660 272576 87712
rect 308312 87660 308364 87712
rect 389180 87660 389232 87712
rect 115940 87592 115992 87644
rect 262864 87592 262916 87644
rect 312544 87592 312596 87644
rect 414020 87592 414072 87644
rect 236000 86436 236052 86488
rect 282736 86436 282788 86488
rect 304816 86436 304868 86488
rect 368480 86436 368532 86488
rect 197360 86368 197412 86420
rect 276296 86368 276348 86420
rect 307760 86368 307812 86420
rect 385040 86368 385092 86420
rect 139400 86300 139452 86352
rect 264244 86300 264296 86352
rect 310888 86300 310940 86352
rect 404360 86300 404412 86352
rect 89720 86232 89772 86284
rect 255964 86232 256016 86284
rect 328000 86232 328052 86284
rect 506480 86232 506532 86284
rect 230480 85076 230532 85128
rect 281816 85076 281868 85128
rect 202880 85008 202932 85060
rect 273996 85008 274048 85060
rect 306472 85008 306524 85060
rect 378140 85008 378192 85060
rect 149060 84940 149112 84992
rect 268384 84940 268436 84992
rect 312176 84940 312228 84992
rect 412640 84940 412692 84992
rect 88340 84872 88392 84924
rect 258264 84872 258316 84924
rect 314752 84872 314804 84924
rect 427820 84872 427872 84924
rect 30380 84804 30432 84856
rect 247684 84804 247736 84856
rect 328552 84804 328604 84856
rect 510620 84804 510672 84856
rect 240140 83716 240192 83768
rect 283196 83716 283248 83768
rect 215300 83648 215352 83700
rect 279332 83648 279384 83700
rect 306932 83648 306984 83700
rect 380900 83648 380952 83700
rect 158720 83580 158772 83632
rect 269948 83580 270000 83632
rect 318064 83580 318116 83632
rect 440332 83580 440384 83632
rect 70400 83512 70452 83564
rect 255044 83512 255096 83564
rect 320364 83512 320416 83564
rect 462412 83512 462464 83564
rect 53840 83444 53892 83496
rect 252560 83444 252612 83496
rect 294420 83444 294472 83496
rect 306380 83444 306432 83496
rect 329012 83444 329064 83496
rect 513380 83444 513432 83496
rect 222200 82288 222252 82340
rect 279608 82288 279660 82340
rect 301780 82288 301832 82340
rect 350540 82288 350592 82340
rect 165620 82220 165672 82272
rect 271052 82220 271104 82272
rect 309140 82220 309192 82272
rect 394700 82220 394752 82272
rect 138020 82152 138072 82204
rect 266452 82152 266504 82204
rect 329564 82152 329616 82204
rect 517612 82152 517664 82204
rect 42800 82084 42852 82136
rect 250628 82084 250680 82136
rect 323952 82084 324004 82136
rect 328460 82084 328512 82136
rect 333060 82084 333112 82136
rect 538220 82084 538272 82136
rect 220820 80860 220872 80912
rect 280344 80860 280396 80912
rect 300124 80860 300176 80912
rect 340972 80860 341024 80912
rect 190460 80792 190512 80844
rect 275192 80792 275244 80844
rect 307484 80792 307536 80844
rect 385132 80792 385184 80844
rect 142160 80724 142212 80776
rect 265624 80724 265676 80776
rect 338948 80724 339000 80776
rect 520280 80724 520332 80776
rect 120080 80656 120132 80708
rect 263324 80656 263376 80708
rect 330300 80656 330352 80708
rect 521660 80656 521712 80708
rect 302240 79500 302292 79552
rect 352012 79500 352064 79552
rect 202972 79432 203024 79484
rect 277676 79432 277728 79484
rect 311348 79432 311400 79484
rect 407120 79432 407172 79484
rect 146300 79364 146352 79416
rect 267740 79364 267792 79416
rect 313280 79364 313332 79416
rect 418160 79364 418212 79416
rect 96620 79296 96672 79348
rect 259460 79296 259512 79348
rect 331772 79296 331824 79348
rect 529940 79296 529992 79348
rect 207020 78140 207072 78192
rect 277952 78140 278004 78192
rect 303252 78140 303304 78192
rect 358820 78140 358872 78192
rect 153200 78072 153252 78124
rect 268844 78072 268896 78124
rect 313004 78072 313056 78124
rect 418252 78072 418304 78124
rect 99380 78004 99432 78056
rect 260012 78004 260064 78056
rect 317052 78004 317104 78056
rect 441620 78004 441672 78056
rect 78680 77936 78732 77988
rect 256516 77936 256568 77988
rect 332324 77936 332376 77988
rect 534080 77936 534132 77988
rect 226340 76712 226392 76764
rect 281172 76712 281224 76764
rect 300492 76712 300544 76764
rect 342260 76712 342312 76764
rect 162860 76644 162912 76696
rect 270500 76644 270552 76696
rect 305460 76644 305512 76696
rect 372620 76644 372672 76696
rect 82820 76576 82872 76628
rect 257252 76576 257304 76628
rect 326344 76576 326396 76628
rect 437480 76576 437532 76628
rect 35900 76508 35952 76560
rect 249340 76508 249392 76560
rect 337476 76508 337528 76560
rect 546500 76508 546552 76560
rect 354404 75828 354456 75880
rect 580172 75828 580224 75880
rect 236092 75352 236144 75404
rect 283012 75352 283064 75404
rect 169852 75284 169904 75336
rect 271144 75284 271196 75336
rect 301596 75284 301648 75336
rect 349160 75284 349212 75336
rect 103520 75216 103572 75268
rect 261024 75216 261076 75268
rect 310980 75216 311032 75268
rect 405740 75216 405792 75268
rect 26240 75148 26292 75200
rect 246396 75148 246448 75200
rect 314108 75148 314160 75200
rect 423680 75148 423732 75200
rect 3332 74468 3384 74520
rect 230020 74468 230072 74520
rect 225052 73924 225104 73976
rect 280804 73924 280856 73976
rect 305000 73924 305052 73976
rect 368572 73924 368624 73976
rect 200120 73856 200172 73908
rect 276848 73856 276900 73908
rect 321560 73856 321612 73908
rect 467932 73856 467984 73908
rect 91100 73788 91152 73840
rect 258632 73788 258684 73840
rect 276020 73788 276072 73840
rect 289452 73788 289504 73840
rect 335084 73788 335136 73840
rect 549904 73788 549956 73840
rect 302700 72632 302752 72684
rect 356060 72632 356112 72684
rect 176660 72564 176712 72616
rect 272892 72564 272944 72616
rect 308772 72564 308824 72616
rect 391940 72564 391992 72616
rect 153292 72496 153344 72548
rect 269304 72496 269356 72548
rect 324412 72496 324464 72548
rect 485780 72496 485832 72548
rect 46940 72428 46992 72480
rect 251180 72428 251232 72480
rect 298836 72428 298888 72480
rect 332600 72428 332652 72480
rect 337384 72428 337436 72480
rect 553400 72428 553452 72480
rect 197452 71136 197504 71188
rect 276388 71136 276440 71188
rect 309692 71136 309744 71188
rect 397460 71136 397512 71188
rect 180800 71068 180852 71120
rect 273536 71068 273588 71120
rect 316500 71068 316552 71120
rect 438860 71068 438912 71120
rect 109040 71000 109092 71052
rect 261668 71000 261720 71052
rect 273260 71000 273312 71052
rect 288992 71000 289044 71052
rect 319628 71000 319680 71052
rect 456892 71000 456944 71052
rect 201500 69776 201552 69828
rect 276940 69776 276992 69828
rect 310244 69776 310296 69828
rect 401600 69776 401652 69828
rect 183560 69708 183612 69760
rect 273628 69708 273680 69760
rect 320180 69708 320232 69760
rect 460940 69708 460992 69760
rect 113180 69640 113232 69692
rect 260104 69640 260156 69692
rect 294972 69640 295024 69692
rect 309140 69640 309192 69692
rect 322756 69640 322808 69692
rect 476120 69640 476172 69692
rect 234620 68484 234672 68536
rect 282460 68484 282512 68536
rect 186320 68416 186372 68468
rect 274916 68416 274968 68468
rect 315212 68416 315264 68468
rect 430580 68416 430632 68468
rect 86960 68348 87012 68400
rect 257804 68348 257856 68400
rect 324780 68348 324832 68400
rect 488540 68348 488592 68400
rect 57980 68280 58032 68332
rect 253020 68280 253072 68332
rect 332784 68280 332836 68332
rect 535460 68280 535512 68332
rect 193220 66988 193272 67040
rect 275652 66988 275704 67040
rect 303988 66988 304040 67040
rect 363052 66988 363104 67040
rect 114560 66920 114612 66972
rect 262496 66920 262548 66972
rect 315764 66920 315816 66972
rect 434812 66920 434864 66972
rect 20720 66852 20772 66904
rect 243636 66852 243688 66904
rect 325884 66852 325936 66904
rect 495440 66852 495492 66904
rect 214012 65628 214064 65680
rect 279148 65628 279200 65680
rect 309508 65628 309560 65680
rect 396080 65628 396132 65680
rect 140780 65560 140832 65612
rect 266820 65560 266872 65612
rect 317420 65560 317472 65612
rect 444380 65560 444432 65612
rect 59360 65492 59412 65544
rect 253388 65492 253440 65544
rect 327540 65492 327592 65544
rect 505100 65492 505152 65544
rect 209780 64268 209832 64320
rect 278412 64268 278464 64320
rect 314476 64268 314528 64320
rect 426440 64268 426492 64320
rect 161480 64200 161532 64252
rect 270316 64200 270368 64252
rect 317972 64200 318024 64252
rect 447140 64200 447192 64252
rect 49700 64132 49752 64184
rect 251732 64132 251784 64184
rect 296812 64132 296864 64184
rect 320180 64132 320232 64184
rect 330852 64132 330904 64184
rect 524420 64132 524472 64184
rect 266452 62976 266504 63028
rect 287796 62976 287848 63028
rect 312268 62908 312320 62960
rect 412732 62908 412784 62960
rect 143540 62840 143592 62892
rect 267372 62840 267424 62892
rect 318524 62840 318576 62892
rect 451280 62840 451332 62892
rect 103612 62772 103664 62824
rect 260564 62772 260616 62824
rect 296260 62772 296312 62824
rect 317420 62772 317472 62824
rect 332692 62772 332744 62824
rect 534172 62772 534224 62824
rect 354312 62024 354364 62076
rect 580172 62024 580224 62076
rect 242900 61548 242952 61600
rect 283932 61548 283984 61600
rect 171140 61480 171192 61532
rect 272064 61480 272116 61532
rect 299480 61480 299532 61532
rect 335360 61480 335412 61532
rect 122840 61412 122892 61464
rect 263876 61412 263928 61464
rect 304356 61412 304408 61464
rect 365720 61412 365772 61464
rect 35164 61344 35216 61396
rect 248880 61344 248932 61396
rect 319260 61344 319312 61396
rect 455420 61344 455472 61396
rect 313372 60120 313424 60172
rect 419540 60120 419592 60172
rect 147680 60052 147732 60104
rect 268016 60052 268068 60104
rect 320732 60052 320784 60104
rect 463700 60052 463752 60104
rect 125600 59984 125652 60036
rect 264428 59984 264480 60036
rect 295708 59984 295760 60036
rect 313280 59984 313332 60036
rect 335820 59984 335872 60036
rect 552664 59984 552716 60036
rect 306564 58760 306616 58812
rect 379520 58760 379572 58812
rect 150440 58692 150492 58744
rect 268476 58692 268528 58744
rect 322020 58692 322072 58744
rect 471980 58692 472032 58744
rect 129740 58624 129792 58676
rect 265072 58624 265124 58676
rect 327172 58624 327224 58676
rect 502340 58624 502392 58676
rect 307116 57332 307168 57384
rect 382280 57332 382332 57384
rect 157340 57264 157392 57316
rect 269580 57264 269632 57316
rect 322572 57264 322624 57316
rect 474740 57264 474792 57316
rect 132500 57196 132552 57248
rect 265164 57196 265216 57248
rect 331036 57196 331088 57248
rect 525800 57196 525852 57248
rect 309324 55972 309376 56024
rect 396172 55972 396224 56024
rect 160100 55904 160152 55956
rect 270132 55904 270184 55956
rect 323124 55904 323176 55956
rect 478880 55904 478932 55956
rect 53932 55836 53984 55888
rect 252284 55836 252336 55888
rect 334348 55836 334400 55888
rect 545120 55836 545172 55888
rect 164240 54544 164292 54596
rect 270776 54544 270828 54596
rect 313740 54544 313792 54596
rect 422300 54544 422352 54596
rect 22100 54476 22152 54528
rect 247408 54476 247460 54528
rect 297180 54476 297232 54528
rect 322940 54476 322992 54528
rect 323676 54476 323728 54528
rect 481640 54476 481692 54528
rect 167000 53116 167052 53168
rect 271236 53116 271288 53168
rect 310520 53116 310572 53168
rect 401692 53116 401744 53168
rect 70492 53048 70544 53100
rect 255504 53048 255556 53100
rect 324320 53048 324372 53100
rect 484492 53048 484544 53100
rect 175372 51756 175424 51808
rect 272616 51756 272668 51808
rect 309876 51756 309928 51808
rect 398840 51756 398892 51808
rect 67640 51688 67692 51740
rect 254676 51688 254728 51740
rect 338856 51688 338908 51740
rect 470600 51688 470652 51740
rect 178040 50396 178092 50448
rect 273076 50396 273128 50448
rect 325332 50396 325384 50448
rect 491300 50396 491352 50448
rect 74540 50328 74592 50380
rect 255872 50328 255924 50380
rect 326068 50328 326120 50380
rect 495532 50328 495584 50380
rect 3240 49648 3292 49700
rect 229928 49648 229980 49700
rect 354220 49648 354272 49700
rect 580172 49648 580224 49700
rect 227720 49036 227772 49088
rect 281356 49036 281408 49088
rect 306012 49036 306064 49088
rect 375380 49036 375432 49088
rect 131120 48968 131172 49020
rect 265256 48968 265308 49020
rect 311716 48968 311768 49020
rect 409880 48968 409932 49020
rect 180892 47608 180944 47660
rect 273720 47608 273772 47660
rect 326436 47608 326488 47660
rect 498200 47608 498252 47660
rect 93860 47540 93912 47592
rect 259092 47540 259144 47592
rect 328828 47540 328880 47592
rect 512000 47540 512052 47592
rect 184940 46248 184992 46300
rect 274180 46248 274232 46300
rect 327080 46248 327132 46300
rect 500960 46248 501012 46300
rect 31760 46180 31812 46232
rect 248604 46180 248656 46232
rect 298468 46180 298520 46232
rect 329840 46180 329892 46232
rect 329932 46180 329984 46232
rect 518900 46180 518952 46232
rect 191932 44888 191984 44940
rect 275100 44888 275152 44940
rect 328092 44888 328144 44940
rect 507860 44888 507912 44940
rect 107660 44820 107712 44872
rect 260932 44820 260984 44872
rect 297916 44820 297968 44872
rect 327080 44820 327132 44872
rect 333796 44820 333848 44872
rect 542360 44820 542412 44872
rect 142252 43460 142304 43512
rect 267004 43460 267056 43512
rect 328644 43460 328696 43512
rect 512092 43460 512144 43512
rect 120172 43392 120224 43444
rect 263784 43392 263836 43444
rect 335452 43392 335504 43444
rect 552020 43392 552072 43444
rect 204260 42100 204312 42152
rect 276664 42100 276716 42152
rect 329196 42100 329248 42152
rect 514760 42100 514812 42152
rect 117320 42032 117372 42084
rect 262956 42032 263008 42084
rect 336004 42032 336056 42084
rect 556252 42032 556304 42084
rect 301228 40808 301280 40860
rect 346492 40808 346544 40860
rect 211160 40740 211212 40792
rect 278596 40740 278648 40792
rect 311164 40740 311216 40792
rect 407212 40740 407264 40792
rect 110420 40672 110472 40724
rect 261852 40672 261904 40724
rect 331404 40672 331456 40724
rect 528560 40672 528612 40724
rect 303436 39448 303488 39500
rect 360200 39448 360252 39500
rect 218060 39380 218112 39432
rect 279700 39380 279752 39432
rect 312820 39380 312872 39432
rect 416780 39380 416832 39432
rect 84200 39312 84252 39364
rect 257528 39312 257580 39364
rect 331956 39312 332008 39364
rect 531320 39312 531372 39364
rect 230572 37952 230624 38004
rect 281908 37952 281960 38004
rect 304540 37952 304592 38004
rect 367100 37952 367152 38004
rect 38660 37884 38712 37936
rect 246304 37884 246356 37936
rect 333612 37884 333664 37936
rect 540980 37884 541032 37936
rect 144920 36592 144972 36644
rect 267556 36592 267608 36644
rect 305092 36592 305144 36644
rect 369860 36592 369912 36644
rect 44180 36524 44232 36576
rect 250812 36524 250864 36576
rect 334164 36524 334216 36576
rect 545212 36524 545264 36576
rect 3332 35844 3384 35896
rect 229836 35844 229888 35896
rect 354128 35844 354180 35896
rect 580172 35844 580224 35896
rect 299020 35232 299072 35284
rect 333980 35232 334032 35284
rect 133880 35164 133932 35216
rect 265808 35164 265860 35216
rect 306196 35164 306248 35216
rect 376760 35164 376812 35216
rect 302332 33872 302384 33924
rect 353300 33872 353352 33924
rect 151820 33804 151872 33856
rect 268660 33804 268712 33856
rect 313924 33804 313976 33856
rect 423772 33804 423824 33856
rect 48320 33736 48372 33788
rect 251456 33736 251508 33788
rect 334716 33736 334768 33788
rect 547880 33736 547932 33788
rect 92572 32444 92624 32496
rect 258724 32444 258776 32496
rect 308404 32444 308456 32496
rect 390652 32444 390704 32496
rect 34520 32376 34572 32428
rect 235264 32376 235316 32428
rect 297364 32376 297416 32428
rect 324320 32376 324372 32428
rect 336372 32376 336424 32428
rect 557540 32376 557592 32428
rect 95240 31084 95292 31136
rect 259276 31084 259328 31136
rect 311532 31084 311584 31136
rect 408500 31084 408552 31136
rect 32404 31016 32456 31068
rect 247868 31016 247920 31068
rect 323308 31016 323360 31068
rect 478972 31016 479024 31068
rect 102140 29656 102192 29708
rect 260380 29656 260432 29708
rect 312636 29656 312688 29708
rect 415400 29656 415452 29708
rect 64880 29588 64932 29640
rect 254124 29588 254176 29640
rect 323860 29588 323912 29640
rect 483020 29588 483072 29640
rect 111800 28296 111852 28348
rect 262036 28296 262088 28348
rect 314292 28296 314344 28348
rect 425060 28296 425112 28348
rect 77300 28228 77352 28280
rect 256332 28228 256384 28280
rect 324964 28228 325016 28280
rect 490012 28228 490064 28280
rect 114652 26936 114704 26988
rect 262680 26936 262732 26988
rect 314844 26936 314896 26988
rect 429292 26936 429344 26988
rect 81532 26868 81584 26920
rect 257160 26868 257212 26920
rect 325516 26868 325568 26920
rect 492680 26868 492732 26920
rect 125692 25576 125744 25628
rect 264336 25576 264388 25628
rect 315396 25576 315448 25628
rect 431960 25576 432012 25628
rect 98092 25508 98144 25560
rect 259552 25508 259604 25560
rect 326620 25508 326672 25560
rect 499580 25508 499632 25560
rect 118700 24148 118752 24200
rect 263140 24148 263192 24200
rect 317604 24148 317656 24200
rect 445852 24148 445904 24200
rect 87052 24080 87104 24132
rect 257344 24080 257396 24132
rect 327724 24080 327776 24132
rect 506572 24080 506624 24132
rect 354036 23400 354088 23452
rect 580172 23400 580224 23452
rect 168380 22788 168432 22840
rect 271420 22788 271472 22840
rect 299572 22788 299624 22840
rect 336832 22788 336884 22840
rect 60740 22720 60792 22772
rect 253572 22720 253624 22772
rect 307300 22720 307352 22772
rect 383660 22720 383712 22772
rect 164332 21428 164384 21480
rect 270960 21428 271012 21480
rect 318156 21428 318208 21480
rect 448520 21428 448572 21480
rect 27620 21360 27672 21412
rect 248052 21360 248104 21412
rect 328276 21360 328328 21412
rect 509240 21360 509292 21412
rect 154580 20000 154632 20052
rect 269212 20000 269264 20052
rect 319812 20000 319864 20052
rect 458180 20000 458232 20052
rect 71780 19932 71832 19984
rect 255412 19932 255464 19984
rect 330484 19932 330536 19984
rect 523040 19932 523092 19984
rect 147772 18640 147824 18692
rect 268292 18640 268344 18692
rect 320916 18640 320968 18692
rect 465080 18640 465132 18692
rect 76012 18572 76064 18624
rect 256056 18572 256108 18624
rect 331588 18572 331640 18624
rect 528652 18572 528704 18624
rect 244280 17348 244332 17400
rect 284116 17348 284168 17400
rect 109132 17280 109184 17332
rect 261576 17280 261628 17332
rect 321652 17280 321704 17332
rect 469220 17280 469272 17332
rect 73160 17212 73212 17264
rect 244924 17212 244976 17264
rect 333244 17212 333296 17264
rect 539692 17212 539744 17264
rect 241704 15920 241756 15972
rect 283380 15920 283432 15972
rect 322204 15920 322256 15972
rect 473544 15920 473596 15972
rect 101496 15852 101548 15904
rect 260196 15852 260248 15904
rect 334900 15852 334952 15904
rect 549720 15852 549772 15904
rect 208584 14492 208636 14544
rect 277860 14492 277912 14544
rect 325056 14492 325108 14544
rect 451372 14492 451424 14544
rect 124680 14424 124732 14476
rect 263692 14424 263744 14476
rect 295156 14424 295208 14476
rect 311256 14424 311308 14476
rect 329380 14424 329432 14476
rect 516600 14424 516652 14476
rect 195336 13132 195388 13184
rect 275836 13132 275888 13184
rect 308956 13132 309008 13184
rect 394056 13132 394108 13184
rect 127992 13064 128044 13116
rect 264612 13064 264664 13116
rect 298284 13064 298336 13116
rect 330024 13064 330076 13116
rect 340144 13064 340196 13116
rect 550732 13064 550784 13116
rect 158904 11772 158956 11824
rect 269764 11772 269816 11824
rect 306748 11772 306800 11824
rect 379612 11772 379664 11824
rect 69480 11704 69532 11756
rect 254860 11704 254912 11756
rect 263784 11704 263836 11756
rect 286324 11704 286376 11756
rect 297732 11704 297784 11756
rect 326712 11704 326764 11756
rect 338764 11704 338816 11756
rect 537576 11704 537628 11756
rect 300216 10956 300268 11008
rect 304172 10956 304224 11008
rect 186504 10344 186556 10396
rect 239404 10344 239456 10396
rect 247408 10344 247460 10396
rect 284668 10344 284720 10396
rect 310060 10344 310112 10396
rect 400680 10344 400732 10396
rect 51816 10276 51868 10328
rect 251916 10276 251968 10328
rect 257160 10276 257212 10328
rect 286140 10276 286192 10328
rect 293316 10276 293368 10328
rect 300216 10276 300268 10328
rect 300676 10276 300728 10328
rect 344376 10276 344428 10328
rect 347044 10276 347096 10328
rect 523132 10276 523184 10328
rect 3424 9596 3476 9648
rect 229744 9596 229796 9648
rect 353944 9596 353996 9648
rect 580172 9596 580224 9648
rect 229560 9528 229612 9580
rect 238024 9528 238076 9580
rect 105912 9120 105964 9172
rect 261484 9120 261536 9172
rect 279240 9120 279292 9172
rect 289176 9120 289228 9172
rect 260472 9052 260524 9104
rect 286692 9052 286744 9104
rect 247224 8984 247276 9036
rect 283656 8984 283708 9036
rect 296720 8984 296772 9036
rect 320088 8984 320140 9036
rect 261576 8916 261628 8968
rect 286876 8916 286928 8968
rect 302884 8916 302936 8968
rect 357624 8916 357676 8968
rect 251640 7692 251692 7744
rect 285220 7692 285272 7744
rect 173256 7624 173308 7676
rect 242164 7624 242216 7676
rect 250536 7624 250588 7676
rect 285036 7624 285088 7676
rect 305644 7624 305696 7676
rect 374184 7624 374236 7676
rect 66168 7556 66220 7608
rect 254400 7556 254452 7608
rect 265992 7556 266044 7608
rect 287152 7556 287204 7608
rect 296444 7556 296496 7608
rect 318984 7556 319036 7608
rect 345664 7556 345716 7608
rect 501144 7556 501196 7608
rect 275928 6876 275980 6928
rect 279516 6876 279568 6928
rect 270408 6400 270460 6452
rect 278044 6400 278096 6452
rect 253848 6332 253900 6384
rect 275284 6332 275336 6384
rect 262680 6264 262732 6316
rect 284944 6264 284996 6316
rect 304448 6264 304500 6316
rect 313464 6264 313516 6316
rect 20904 6196 20956 6248
rect 245752 6196 245804 6248
rect 258264 6196 258316 6248
rect 286416 6196 286468 6248
rect 294604 6196 294656 6248
rect 307944 6196 307996 6248
rect 342904 6196 342956 6248
rect 487896 6196 487948 6248
rect 19800 6128 19852 6180
rect 245660 6128 245712 6180
rect 252744 6128 252796 6180
rect 285404 6128 285456 6180
rect 285864 6128 285916 6180
rect 290924 6128 290976 6180
rect 295892 6128 295944 6180
rect 315672 6128 315724 6180
rect 332140 6128 332192 6180
rect 533160 6128 533212 6180
rect 280344 5516 280396 5568
rect 289084 5516 289136 5568
rect 272616 5108 272668 5160
rect 282276 5108 282328 5160
rect 269304 5040 269356 5092
rect 288164 5040 288216 5092
rect 256056 4972 256108 5024
rect 273904 4972 273956 5024
rect 136824 4904 136876 4956
rect 254952 4904 255004 4956
rect 283564 4904 283616 4956
rect 293684 4904 293736 4956
rect 302424 4904 302476 4956
rect 243544 4836 243596 4888
rect 249432 4836 249484 4888
rect 282184 4836 282236 4888
rect 295340 4836 295392 4888
rect 312360 4836 312412 4888
rect 341524 4836 341576 4888
rect 474648 4836 474700 4888
rect 475384 4836 475436 4888
rect 497832 4836 497884 4888
rect 86040 4768 86092 4820
rect 257620 4768 257672 4820
rect 259368 4768 259420 4820
rect 279424 4768 279476 4820
rect 296076 4768 296128 4820
rect 316776 4768 316828 4820
rect 323768 4768 323820 4820
rect 335544 4768 335596 4820
rect 336556 4768 336608 4820
rect 559656 4768 559708 4820
rect 301688 4496 301740 4548
rect 309048 4496 309100 4548
rect 282552 4428 282604 4480
rect 287704 4428 287756 4480
rect 293132 4360 293184 4412
rect 299112 4360 299164 4412
rect 70492 4156 70544 4208
rect 71688 4156 71740 4208
rect 87052 4156 87104 4208
rect 88248 4156 88300 4208
rect 114652 4156 114704 4208
rect 115848 4156 115900 4208
rect 120172 4156 120224 4208
rect 121368 4156 121420 4208
rect 147772 4156 147824 4208
rect 148968 4156 149020 4208
rect 153292 4156 153344 4208
rect 154488 4156 154540 4208
rect 164332 4156 164384 4208
rect 165528 4156 165580 4208
rect 169852 4156 169904 4208
rect 171048 4156 171100 4208
rect 180892 4156 180944 4208
rect 182088 4156 182140 4208
rect 197452 4156 197504 4208
rect 198648 4156 198700 4208
rect 202972 4156 203024 4208
rect 204168 4156 204220 4208
rect 214012 4156 214064 4208
rect 215208 4156 215260 4208
rect 230572 4156 230624 4208
rect 231768 4156 231820 4208
rect 236092 4156 236144 4208
rect 237288 4156 237340 4208
rect 301504 4156 301556 4208
rect 303528 4156 303580 4208
rect 304264 4156 304316 4208
rect 305736 4156 305788 4208
rect 320824 4156 320876 4208
rect 322296 4156 322348 4208
rect 323584 4156 323636 4208
rect 325608 4156 325660 4208
rect 346492 4156 346544 4208
rect 347688 4156 347740 4208
rect 352012 4156 352064 4208
rect 353208 4156 353260 4208
rect 363052 4156 363104 4208
rect 364248 4156 364300 4208
rect 368572 4156 368624 4208
rect 369768 4156 369820 4208
rect 379612 4156 379664 4208
rect 380808 4156 380860 4208
rect 401692 4156 401744 4208
rect 402888 4156 402940 4208
rect 412732 4156 412784 4208
rect 413928 4156 413980 4208
rect 59544 4088 59596 4140
rect 253204 4088 253256 4140
rect 292948 4088 293000 4140
rect 298008 4088 298060 4140
rect 316684 4088 316736 4140
rect 440424 4088 440476 4140
rect 56232 4020 56284 4072
rect 252652 4020 252704 4072
rect 317236 4020 317288 4072
rect 443736 4020 443788 4072
rect 451372 4020 451424 4072
rect 452568 4020 452620 4072
rect 52920 3952 52972 4004
rect 252100 3952 252152 4004
rect 284760 3952 284812 4004
rect 290740 3952 290792 4004
rect 317788 3952 317840 4004
rect 447048 3952 447100 4004
rect 25320 3884 25372 3936
rect 28264 3884 28316 3936
rect 49608 3884 49660 3936
rect 251548 3884 251600 3936
rect 286968 3884 287020 3936
rect 291384 3884 291436 3936
rect 292764 3884 292816 3936
rect 296904 3884 296956 3936
rect 318340 3884 318392 3936
rect 450360 3884 450412 3936
rect 46296 3816 46348 3868
rect 250996 3816 251048 3868
rect 283656 3816 283708 3868
rect 290556 3816 290608 3868
rect 318892 3816 318944 3868
rect 453672 3952 453724 4004
rect 42984 3748 43036 3800
rect 250444 3748 250496 3800
rect 281448 3748 281500 3800
rect 290188 3748 290240 3800
rect 319444 3748 319496 3800
rect 456984 3748 457036 3800
rect 41880 3680 41932 3732
rect 250260 3680 250312 3732
rect 278136 3680 278188 3732
rect 289636 3680 289688 3732
rect 319996 3680 320048 3732
rect 460296 3680 460348 3732
rect 38568 3612 38620 3664
rect 33048 3544 33100 3596
rect 35164 3544 35216 3596
rect 42800 3544 42852 3596
rect 44088 3544 44140 3596
rect 44272 3612 44324 3664
rect 249524 3612 249576 3664
rect 274824 3612 274876 3664
rect 288624 3612 288676 3664
rect 292396 3612 292448 3664
rect 294696 3612 294748 3664
rect 320548 3612 320600 3664
rect 463608 3612 463660 3664
rect 467932 3612 467984 3664
rect 469128 3612 469180 3664
rect 478972 3612 479024 3664
rect 480168 3612 480220 3664
rect 484492 3612 484544 3664
rect 485688 3612 485740 3664
rect 495532 3612 495584 3664
rect 496728 3612 496780 3664
rect 523132 3612 523184 3664
rect 524328 3612 524380 3664
rect 528652 3612 528704 3664
rect 529848 3612 529900 3664
rect 534172 3612 534224 3664
rect 535368 3612 535420 3664
rect 552664 3612 552716 3664
rect 555240 3612 555292 3664
rect 249984 3544 250036 3596
rect 271512 3544 271564 3596
rect 288900 3544 288952 3596
rect 292212 3544 292264 3596
rect 293592 3544 293644 3596
rect 336924 3544 336976 3596
rect 562968 3544 563020 3596
rect 34152 3476 34204 3528
rect 248972 3476 249024 3528
rect 268200 3476 268252 3528
rect 287980 3476 288032 3528
rect 288072 3476 288124 3528
rect 291476 3476 291528 3528
rect 313280 3476 313332 3528
rect 314568 3476 314620 3528
rect 321284 3476 321336 3528
rect 466920 3476 466972 3528
rect 489920 3476 489972 3528
rect 491208 3476 491260 3528
rect 500960 3476 501012 3528
rect 502248 3476 502300 3528
rect 506480 3476 506532 3528
rect 507768 3476 507820 3528
rect 512000 3476 512052 3528
rect 513288 3476 513340 3528
rect 517520 3476 517572 3528
rect 518808 3476 518860 3528
rect 549904 3476 549956 3528
rect 550824 3476 550876 3528
rect 29736 3408 29788 3460
rect 241428 3408 241480 3460
rect 241520 3408 241572 3460
rect 242808 3408 242860 3460
rect 264888 3408 264940 3460
rect 287520 3408 287572 3460
rect 290280 3408 290332 3460
rect 291752 3408 291804 3460
rect 293500 3408 293552 3460
rect 301320 3408 301372 3460
rect 340880 3408 340932 3460
rect 342168 3408 342220 3460
rect 342260 3408 342312 3460
rect 561864 3408 561916 3460
rect 37464 3340 37516 3392
rect 44272 3340 44324 3392
rect 53840 3340 53892 3392
rect 55128 3340 55180 3392
rect 59360 3340 59412 3392
rect 60648 3340 60700 3392
rect 62856 3340 62908 3392
rect 253756 3340 253808 3392
rect 292580 3340 292632 3392
rect 295800 3340 295852 3392
rect 316132 3340 316184 3392
rect 75920 3272 75972 3324
rect 77208 3272 77260 3324
rect 81440 3272 81492 3324
rect 82728 3272 82780 3324
rect 92480 3272 92532 3324
rect 93768 3272 93820 3324
rect 98000 3272 98052 3324
rect 99288 3272 99340 3324
rect 103520 3272 103572 3324
rect 104808 3272 104860 3324
rect 109040 3272 109092 3324
rect 110328 3272 110380 3324
rect 125600 3272 125652 3324
rect 126888 3272 126940 3324
rect 132408 3272 132460 3324
rect 265532 3272 265584 3324
rect 315580 3272 315632 3324
rect 433800 3272 433852 3324
rect 434720 3340 434772 3392
rect 436008 3340 436060 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 456892 3340 456944 3392
rect 458088 3340 458140 3392
rect 550732 3340 550784 3392
rect 551928 3340 551980 3392
rect 437112 3272 437164 3324
rect 135720 3204 135772 3256
rect 265900 3204 265952 3256
rect 315028 3204 315080 3256
rect 142160 3136 142212 3188
rect 143448 3136 143500 3188
rect 158720 3136 158772 3188
rect 160008 3136 160060 3188
rect 175280 3136 175332 3188
rect 176568 3136 176620 3188
rect 186320 3136 186372 3188
rect 187608 3136 187660 3188
rect 191840 3136 191892 3188
rect 193128 3136 193180 3188
rect 208400 3136 208452 3188
rect 209688 3136 209740 3188
rect 219440 3136 219492 3188
rect 220728 3136 220780 3188
rect 224960 3136 225012 3188
rect 226248 3136 226300 3188
rect 241428 3136 241480 3188
rect 248236 3136 248288 3188
rect 289176 3136 289228 3188
rect 291568 3136 291620 3188
rect 336740 3136 336792 3188
rect 342260 3136 342312 3188
rect 357440 3136 357492 3188
rect 358728 3136 358780 3188
rect 374000 3136 374052 3188
rect 375288 3136 375340 3188
rect 385040 3136 385092 3188
rect 386328 3136 386380 3188
rect 390560 3136 390612 3188
rect 391848 3136 391900 3188
rect 396080 3136 396132 3188
rect 397368 3136 397420 3188
rect 407120 3136 407172 3188
rect 408408 3136 408460 3188
rect 418160 3204 418212 3256
rect 419448 3204 419500 3256
rect 423680 3204 423732 3256
rect 424968 3204 425020 3256
rect 430488 3136 430540 3188
rect 27528 3000 27580 3052
rect 32404 3000 32456 3052
rect 136640 2728 136692 2780
rect 137928 2728 137980 2780
rect 335360 2592 335412 2644
rect 336648 2592 336700 2644
rect 329840 2388 329892 2440
rect 331128 2388 331180 2440
rect 20720 2320 20772 2372
rect 22008 2320 22060 2372
rect 539600 1232 539652 1284
rect 540888 1232 540940 1284
rect 545120 1232 545172 1284
rect 546408 1232 546460 1284
rect 556160 1232 556212 1284
rect 557448 1232 557500 1284
<< metal2 >>
rect 8546 703520 8658 704960
rect 24738 703520 24850 704960
rect 40930 703520 41042 704960
rect 57122 703520 57234 704960
rect 73314 703520 73426 704960
rect 89506 703520 89618 704960
rect 105698 703520 105810 704960
rect 121890 703520 122002 704960
rect 138082 703520 138194 704960
rect 154274 703520 154386 704960
rect 170466 703520 170578 704960
rect 186658 703520 186770 704960
rect 202850 703520 202962 704960
rect 219042 703520 219154 704960
rect 235234 703520 235346 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300002 703520 300114 704960
rect 316194 703520 316306 704960
rect 332386 703520 332498 704960
rect 348578 703520 348690 704960
rect 364770 703520 364882 704960
rect 380962 703520 381074 704960
rect 397154 703520 397266 704960
rect 413346 703520 413458 704960
rect 429538 703520 429650 704960
rect 445730 703520 445842 704960
rect 461922 703520 462034 704960
rect 478114 703520 478226 704960
rect 494306 703520 494418 704960
rect 510498 703520 510610 704960
rect 526690 703520 526802 704960
rect 542882 703520 542994 704960
rect 559074 703520 559186 704960
rect 575266 703520 575378 704960
rect 8588 702434 8616 703520
rect 8312 702406 8616 702434
rect 2778 681456 2834 681465
rect 2778 681391 2834 681400
rect 2792 680610 2820 681391
rect 2780 680604 2832 680610
rect 2780 680546 2832 680552
rect 4804 680604 4856 680610
rect 4804 680546 4856 680552
rect 3422 668536 3478 668545
rect 3422 668471 3478 668480
rect 3330 616856 3386 616865
rect 3330 616791 3386 616800
rect 3344 615534 3372 616791
rect 3332 615528 3384 615534
rect 3332 615470 3384 615476
rect 3330 603936 3386 603945
rect 3330 603871 3386 603880
rect 3344 603158 3372 603871
rect 3332 603152 3384 603158
rect 3332 603094 3384 603100
rect 3330 578096 3386 578105
rect 3330 578031 3386 578040
rect 3344 576910 3372 578031
rect 3332 576904 3384 576910
rect 3332 576846 3384 576852
rect 3330 526416 3386 526425
rect 3330 526351 3386 526360
rect 3344 525842 3372 526351
rect 3332 525836 3384 525842
rect 3332 525778 3384 525784
rect 3330 513496 3386 513505
rect 3330 513431 3386 513440
rect 3344 513398 3372 513431
rect 3332 513392 3384 513398
rect 3332 513334 3384 513340
rect 2962 500576 3018 500585
rect 2962 500511 3018 500520
rect 2976 499594 3004 500511
rect 2964 499588 3016 499594
rect 2964 499530 3016 499536
rect 3238 474736 3294 474745
rect 3238 474671 3294 474680
rect 3252 474094 3280 474671
rect 3240 474088 3292 474094
rect 3240 474030 3292 474036
rect 2962 423056 3018 423065
rect 2962 422991 3018 423000
rect 2976 422346 3004 422991
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3330 410136 3386 410145
rect 3330 410071 3386 410080
rect 3344 409902 3372 410071
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 2962 397216 3018 397225
rect 2962 397151 3018 397160
rect 2976 396098 3004 397151
rect 2964 396092 3016 396098
rect 2964 396034 3016 396040
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 319696 3386 319705
rect 3330 319631 3386 319640
rect 3344 318850 3372 319631
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3330 306776 3386 306785
rect 3330 306711 3386 306720
rect 3344 306406 3372 306711
rect 3332 306400 3384 306406
rect 3332 306342 3384 306348
rect 3330 293856 3386 293865
rect 3330 293791 3386 293800
rect 3344 292602 3372 293791
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3330 268016 3386 268025
rect 3330 267951 3386 267960
rect 3344 267782 3372 267951
rect 3332 267776 3384 267782
rect 3332 267718 3384 267724
rect 3436 255270 3464 668471
rect 3514 655616 3570 655625
rect 3514 655551 3570 655560
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3330 255096 3386 255105
rect 3330 255031 3386 255040
rect 3344 162858 3372 255031
rect 3528 251190 3556 655551
rect 3606 629776 3662 629785
rect 3606 629711 3662 629720
rect 3620 629338 3648 629711
rect 3608 629332 3660 629338
rect 3608 629274 3660 629280
rect 3606 565176 3662 565185
rect 3606 565111 3662 565120
rect 3516 251184 3568 251190
rect 3516 251126 3568 251132
rect 3422 242176 3478 242185
rect 3422 242111 3478 242120
rect 3332 162852 3384 162858
rect 3332 162794 3384 162800
rect 3436 160070 3464 242111
rect 3620 231810 3648 565111
rect 3698 552256 3754 552265
rect 3698 552191 3754 552200
rect 3608 231804 3660 231810
rect 3608 231746 3660 231752
rect 3712 227730 3740 552191
rect 3790 461816 3846 461825
rect 3790 461751 3846 461760
rect 3700 227724 3752 227730
rect 3700 227666 3752 227672
rect 3514 216336 3570 216345
rect 3514 216271 3570 216280
rect 3424 160064 3476 160070
rect 3424 160006 3476 160012
rect 3528 155922 3556 216271
rect 3804 209778 3832 461751
rect 3882 448896 3938 448905
rect 3882 448831 3938 448840
rect 3792 209772 3844 209778
rect 3792 209714 3844 209720
rect 3896 205630 3924 448831
rect 3974 358456 4030 358465
rect 3974 358391 4030 358400
rect 3884 205624 3936 205630
rect 3884 205566 3936 205572
rect 3606 203416 3662 203425
rect 3606 203351 3662 203360
rect 3516 155916 3568 155922
rect 3516 155858 3568 155864
rect 3620 151774 3648 203351
rect 3698 190496 3754 190505
rect 3698 190431 3754 190440
rect 3608 151768 3660 151774
rect 3422 151736 3478 151745
rect 3608 151710 3660 151716
rect 3422 151671 3478 151680
rect 3436 140758 3464 151671
rect 3712 147626 3740 190431
rect 3988 186318 4016 358391
rect 4066 345536 4122 345545
rect 4066 345471 4122 345480
rect 3976 186312 4028 186318
rect 3976 186254 4028 186260
rect 4080 182170 4108 345471
rect 4816 258058 4844 680546
rect 7564 576904 7616 576910
rect 7564 576846 7616 576852
rect 4804 258052 4856 258058
rect 4804 257994 4856 258000
rect 7576 235958 7604 576846
rect 8312 262886 8340 702406
rect 24780 697610 24808 703520
rect 40972 702434 41000 703520
rect 40052 702406 41000 702434
rect 23480 697604 23532 697610
rect 23480 697546 23532 697552
rect 24768 697604 24820 697610
rect 24768 697546 24820 697552
rect 22744 615528 22796 615534
rect 22744 615470 22796 615476
rect 14464 603152 14516 603158
rect 14464 603094 14516 603100
rect 8944 474088 8996 474094
rect 8944 474030 8996 474036
rect 8300 262880 8352 262886
rect 8300 262822 8352 262828
rect 7564 235952 7616 235958
rect 7564 235894 7616 235900
rect 8956 212498 8984 474030
rect 10324 371272 10376 371278
rect 10324 371214 10376 371220
rect 8944 212492 8996 212498
rect 8944 212434 8996 212440
rect 10336 190466 10364 371214
rect 13084 267776 13136 267782
rect 13084 267718 13136 267724
rect 10324 190460 10376 190466
rect 10324 190402 10376 190408
rect 4068 182164 4120 182170
rect 4068 182106 4120 182112
rect 13096 167006 13124 267718
rect 14476 240106 14504 603094
rect 17224 499588 17276 499594
rect 17224 499530 17276 499536
rect 14464 240100 14516 240106
rect 14464 240042 14516 240048
rect 17236 216646 17264 499530
rect 18604 396092 18656 396098
rect 18604 396034 18656 396040
rect 17224 216640 17276 216646
rect 17224 216582 17276 216588
rect 18616 193186 18644 396034
rect 21364 292596 21416 292602
rect 21364 292538 21416 292544
rect 18604 193180 18656 193186
rect 18604 193122 18656 193128
rect 21376 171086 21404 292538
rect 22756 242894 22784 615470
rect 23492 262954 23520 697546
rect 35164 629332 35216 629338
rect 35164 629274 35216 629280
rect 25504 513392 25556 513398
rect 25504 513334 25556 513340
rect 23480 262948 23532 262954
rect 23480 262890 23532 262896
rect 22744 242888 22796 242894
rect 22744 242830 22796 242836
rect 25516 220794 25544 513334
rect 26884 409896 26936 409902
rect 26884 409838 26936 409844
rect 25504 220788 25556 220794
rect 25504 220730 25556 220736
rect 26896 197334 26924 409838
rect 28264 306400 28316 306406
rect 28264 306342 28316 306348
rect 26884 197328 26936 197334
rect 26884 197270 26936 197276
rect 28276 175234 28304 306342
rect 35176 247042 35204 629274
rect 40052 263022 40080 702406
rect 73356 683114 73384 703520
rect 89548 703050 89576 703520
rect 88340 703044 88392 703050
rect 88340 702986 88392 702992
rect 89536 703044 89588 703050
rect 89536 702986 89588 702992
rect 73172 683086 73384 683114
rect 61384 525836 61436 525842
rect 61384 525778 61436 525784
rect 40040 263016 40092 263022
rect 40040 262958 40092 262964
rect 35164 247036 35216 247042
rect 35164 246978 35216 246984
rect 61396 224942 61424 525778
rect 73172 263090 73200 683086
rect 88352 263158 88380 702986
rect 105740 702434 105768 703520
rect 104912 702406 105768 702434
rect 104912 263226 104940 702406
rect 138124 683114 138152 703520
rect 154316 702434 154344 703520
rect 170508 702434 170536 703520
rect 138032 683086 138152 683114
rect 153212 702406 154344 702434
rect 169772 702406 170536 702434
rect 138032 263294 138060 683086
rect 153212 263362 153240 702406
rect 169772 263430 169800 702406
rect 180064 422340 180116 422346
rect 180064 422282 180116 422288
rect 169760 263424 169812 263430
rect 169760 263366 169812 263372
rect 153200 263356 153252 263362
rect 153200 263298 153252 263304
rect 138020 263288 138072 263294
rect 138020 263230 138072 263236
rect 104900 263220 104952 263226
rect 104900 263162 104952 263168
rect 88340 263152 88392 263158
rect 88340 263094 88392 263100
rect 73160 263084 73212 263090
rect 73160 263026 73212 263032
rect 61384 224936 61436 224942
rect 61384 224878 61436 224884
rect 180076 201482 180104 422282
rect 202892 263498 202920 703520
rect 219084 702434 219112 703520
rect 235276 702434 235304 703520
rect 218072 702406 219112 702434
rect 234632 702406 235304 702434
rect 218072 263566 218100 702406
rect 224224 318844 224276 318850
rect 224224 318786 224276 318792
rect 218060 263560 218112 263566
rect 218060 263502 218112 263508
rect 202880 263492 202932 263498
rect 202880 263434 202932 263440
rect 180064 201476 180116 201482
rect 180064 201418 180116 201424
rect 224236 178022 224264 318786
rect 234632 262886 234660 702406
rect 267660 700330 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 279424 700324 279476 700330
rect 279424 700266 279476 700272
rect 278688 263560 278740 263566
rect 278688 263502 278740 263508
rect 274272 263492 274324 263498
rect 274272 263434 274324 263440
rect 269856 263424 269908 263430
rect 269856 263366 269908 263372
rect 265440 263356 265492 263362
rect 265440 263298 265492 263304
rect 261024 263288 261076 263294
rect 261024 263230 261076 263236
rect 256608 263220 256660 263226
rect 256608 263162 256660 263168
rect 252192 263152 252244 263158
rect 252192 263094 252244 263100
rect 247776 263084 247828 263090
rect 247776 263026 247828 263032
rect 243360 263016 243412 263022
rect 243360 262958 243412 262964
rect 238944 262948 238996 262954
rect 238944 262890 238996 262896
rect 234528 262880 234580 262886
rect 234528 262822 234580 262828
rect 234620 262880 234672 262886
rect 234620 262822 234672 262828
rect 234540 259964 234568 262822
rect 238956 259964 238984 262890
rect 243372 259964 243400 262958
rect 247788 259964 247816 263026
rect 252204 259964 252232 263094
rect 256620 259964 256648 263162
rect 261036 259964 261064 263230
rect 265452 259964 265480 263298
rect 269868 259964 269896 263366
rect 274284 259964 274312 263434
rect 278700 259964 278728 263502
rect 279436 262954 279464 700266
rect 282932 263022 282960 702406
rect 300044 700534 300072 703520
rect 309140 700936 309192 700942
rect 309140 700878 309192 700884
rect 295340 700528 295392 700534
rect 295340 700470 295392 700476
rect 300032 700528 300084 700534
rect 300032 700470 300084 700476
rect 295352 267734 295380 700470
rect 299480 700392 299532 700398
rect 299480 700334 299532 700340
rect 299492 267734 299520 700334
rect 305000 700324 305052 700330
rect 305000 700266 305052 700272
rect 295352 267706 296024 267734
rect 299492 267706 300440 267734
rect 282920 263016 282972 263022
rect 282920 262958 282972 262964
rect 291936 263016 291988 263022
rect 291936 262958 291988 262964
rect 279424 262948 279476 262954
rect 279424 262890 279476 262896
rect 287520 262948 287572 262954
rect 287520 262890 287572 262896
rect 283104 262880 283156 262886
rect 283104 262822 283156 262828
rect 283116 259964 283144 262822
rect 287532 259964 287560 262890
rect 291948 259964 291976 262958
rect 295996 259978 296024 267706
rect 300412 259978 300440 267706
rect 305012 259978 305040 700266
rect 309152 267734 309180 700878
rect 313280 700868 313332 700874
rect 313280 700810 313332 700816
rect 313292 267734 313320 700810
rect 317420 700800 317472 700806
rect 317420 700742 317472 700748
rect 317432 267734 317460 700742
rect 321560 700732 321612 700738
rect 321560 700674 321612 700680
rect 321572 267734 321600 700674
rect 327080 700664 327132 700670
rect 327080 700606 327132 700612
rect 309152 267706 309272 267734
rect 313292 267706 313688 267734
rect 317432 267706 318104 267734
rect 321572 267706 322520 267734
rect 309244 259978 309272 267706
rect 313660 259978 313688 267706
rect 318076 259978 318104 267706
rect 322492 259978 322520 267706
rect 327092 259978 327120 700606
rect 331312 700596 331364 700602
rect 331312 700538 331364 700544
rect 331324 259978 331352 700538
rect 332428 700398 332456 703520
rect 335360 700528 335412 700534
rect 335360 700470 335412 700476
rect 332416 700392 332468 700398
rect 332416 700334 332468 700340
rect 335372 267734 335400 700470
rect 339500 700460 339552 700466
rect 339500 700402 339552 700408
rect 339512 267734 339540 700402
rect 343640 700392 343692 700398
rect 343640 700334 343692 700340
rect 343652 267734 343680 700334
rect 348620 700330 348648 703520
rect 364812 700942 364840 703520
rect 364800 700936 364852 700942
rect 364800 700878 364852 700884
rect 397196 700874 397224 703520
rect 397184 700868 397236 700874
rect 397184 700810 397236 700816
rect 413388 700806 413416 703520
rect 413376 700800 413428 700806
rect 413376 700742 413428 700748
rect 429580 700738 429608 703520
rect 429568 700732 429620 700738
rect 429568 700674 429620 700680
rect 461964 700670 461992 703520
rect 461952 700664 462004 700670
rect 461952 700606 462004 700612
rect 478156 700602 478184 703520
rect 478144 700596 478196 700602
rect 478144 700538 478196 700544
rect 494348 700534 494376 703520
rect 494336 700528 494388 700534
rect 494336 700470 494388 700476
rect 526732 700466 526760 703520
rect 526720 700460 526772 700466
rect 526720 700402 526772 700408
rect 542924 700398 542952 703520
rect 542912 700392 542964 700398
rect 542912 700334 542964 700340
rect 559116 700330 559144 703520
rect 348608 700324 348660 700330
rect 348608 700266 348660 700272
rect 349160 700324 349212 700330
rect 349160 700266 349212 700272
rect 559104 700324 559156 700330
rect 559104 700266 559156 700272
rect 335372 267706 335768 267734
rect 339512 267706 340184 267734
rect 343652 267706 344600 267734
rect 335740 259978 335768 267706
rect 340156 259978 340184 267706
rect 344572 259978 344600 267706
rect 349172 259978 349200 700266
rect 580262 694920 580318 694929
rect 580262 694855 580318 694864
rect 580170 681728 580226 681737
rect 580170 681663 580226 681672
rect 580184 680406 580212 681663
rect 353944 680400 353996 680406
rect 353944 680342 353996 680348
rect 580172 680400 580224 680406
rect 580172 680342 580224 680348
rect 295996 259950 296378 259978
rect 300412 259950 300794 259978
rect 305012 259950 305210 259978
rect 309244 259950 309626 259978
rect 313660 259950 314042 259978
rect 318076 259950 318458 259978
rect 322492 259950 322874 259978
rect 327092 259950 327290 259978
rect 331324 259950 331706 259978
rect 335740 259950 336122 259978
rect 340156 259950 340538 259978
rect 344572 259950 344954 259978
rect 349172 259950 349370 259978
rect 230388 258052 230440 258058
rect 230388 257994 230440 258000
rect 353300 258052 353352 258058
rect 353300 257994 353352 258000
rect 230400 257961 230428 257994
rect 230386 257952 230442 257961
rect 230386 257887 230442 257896
rect 353312 257689 353340 257994
rect 353298 257680 353354 257689
rect 353298 257615 353354 257624
rect 230388 255264 230440 255270
rect 230388 255206 230440 255212
rect 230400 254153 230428 255206
rect 353956 254153 353984 680342
rect 580170 668536 580226 668545
rect 580170 668471 580226 668480
rect 580184 667962 580212 668471
rect 360844 667956 360896 667962
rect 360844 667898 360896 667904
rect 580172 667956 580224 667962
rect 580172 667898 580224 667904
rect 359464 561740 359516 561746
rect 359464 561682 359516 561688
rect 356704 509312 356756 509318
rect 356704 509254 356756 509260
rect 355324 456816 355376 456822
rect 355324 456758 355376 456764
rect 354036 364404 354088 364410
rect 354036 364346 354088 364352
rect 230386 254144 230442 254153
rect 230386 254079 230442 254088
rect 353942 254144 353998 254153
rect 353942 254079 353998 254088
rect 230388 251184 230440 251190
rect 230388 251126 230440 251132
rect 353300 251184 353352 251190
rect 353300 251126 353352 251132
rect 230400 250345 230428 251126
rect 353312 250617 353340 251126
rect 353298 250608 353354 250617
rect 353298 250543 353354 250552
rect 230386 250336 230442 250345
rect 230386 250271 230442 250280
rect 353300 248396 353352 248402
rect 353300 248338 353352 248344
rect 353312 247081 353340 248338
rect 353298 247072 353354 247081
rect 229652 247036 229704 247042
rect 353298 247007 353354 247016
rect 229652 246978 229704 246984
rect 229664 246537 229692 246978
rect 229650 246528 229706 246537
rect 229650 246463 229706 246472
rect 353300 244248 353352 244254
rect 353300 244190 353352 244196
rect 353312 243545 353340 244190
rect 353298 243536 353354 243545
rect 353298 243471 353354 243480
rect 229284 242888 229336 242894
rect 229284 242830 229336 242836
rect 229296 242729 229324 242830
rect 229282 242720 229338 242729
rect 229282 242655 229338 242664
rect 230020 240100 230072 240106
rect 230020 240042 230072 240048
rect 353300 240100 353352 240106
rect 353300 240042 353352 240048
rect 230032 238921 230060 240042
rect 353312 240009 353340 240042
rect 353298 240000 353354 240009
rect 353298 239935 353354 239944
rect 230018 238912 230074 238921
rect 230018 238847 230074 238856
rect 353300 237380 353352 237386
rect 353300 237322 353352 237328
rect 353312 236473 353340 237322
rect 353298 236464 353354 236473
rect 353298 236399 353354 236408
rect 230204 235952 230256 235958
rect 230204 235894 230256 235900
rect 230216 235113 230244 235894
rect 230202 235104 230258 235113
rect 230202 235039 230258 235048
rect 353300 233232 353352 233238
rect 353300 233174 353352 233180
rect 353312 232937 353340 233174
rect 353298 232928 353354 232937
rect 353298 232863 353354 232872
rect 230388 231804 230440 231810
rect 230388 231746 230440 231752
rect 230400 231305 230428 231746
rect 230386 231296 230442 231305
rect 230386 231231 230442 231240
rect 353300 230444 353352 230450
rect 353300 230386 353352 230392
rect 353312 229401 353340 230386
rect 353298 229392 353354 229401
rect 353298 229327 353354 229336
rect 230388 227724 230440 227730
rect 230388 227666 230440 227672
rect 230400 227497 230428 227666
rect 230386 227488 230442 227497
rect 230386 227423 230442 227432
rect 353300 226296 353352 226302
rect 353300 226238 353352 226244
rect 353312 225865 353340 226238
rect 353298 225856 353354 225865
rect 353298 225791 353354 225800
rect 229652 224936 229704 224942
rect 229652 224878 229704 224884
rect 229664 223689 229692 224878
rect 229650 223680 229706 223689
rect 229650 223615 229706 223624
rect 353300 223576 353352 223582
rect 353300 223518 353352 223524
rect 353312 222329 353340 223518
rect 353298 222320 353354 222329
rect 353298 222255 353354 222264
rect 230388 220788 230440 220794
rect 230388 220730 230440 220736
rect 230400 219881 230428 220730
rect 230386 219872 230442 219881
rect 230386 219807 230442 219816
rect 353944 219496 353996 219502
rect 353944 219438 353996 219444
rect 353300 219428 353352 219434
rect 353300 219370 353352 219376
rect 353312 218793 353340 219370
rect 353298 218784 353354 218793
rect 353298 218719 353354 218728
rect 230388 216640 230440 216646
rect 230388 216582 230440 216588
rect 230400 216073 230428 216582
rect 230386 216064 230442 216073
rect 230386 215999 230442 216008
rect 353300 215280 353352 215286
rect 353298 215248 353300 215257
rect 353352 215248 353354 215257
rect 353298 215183 353354 215192
rect 230388 212492 230440 212498
rect 230388 212434 230440 212440
rect 353300 212492 353352 212498
rect 353300 212434 353352 212440
rect 230400 212265 230428 212434
rect 230386 212256 230442 212265
rect 230386 212191 230442 212200
rect 353312 211721 353340 212434
rect 353298 211712 353354 211721
rect 353298 211647 353354 211656
rect 229652 209772 229704 209778
rect 229652 209714 229704 209720
rect 229664 208457 229692 209714
rect 229650 208448 229706 208457
rect 229650 208383 229706 208392
rect 353300 208208 353352 208214
rect 353298 208176 353300 208185
rect 353352 208176 353354 208185
rect 353298 208111 353354 208120
rect 229468 205624 229520 205630
rect 229468 205566 229520 205572
rect 353300 205624 353352 205630
rect 353300 205566 353352 205572
rect 229480 204649 229508 205566
rect 353312 204649 353340 205566
rect 229466 204640 229522 204649
rect 229466 204575 229522 204584
rect 353298 204640 353354 204649
rect 353298 204575 353354 204584
rect 230388 201476 230440 201482
rect 230388 201418 230440 201424
rect 353300 201476 353352 201482
rect 353300 201418 353352 201424
rect 230400 200841 230428 201418
rect 353312 201113 353340 201418
rect 353298 201104 353354 201113
rect 353298 201039 353354 201048
rect 230386 200832 230442 200841
rect 230386 200767 230442 200776
rect 353300 198688 353352 198694
rect 353300 198630 353352 198636
rect 353312 197577 353340 198630
rect 353298 197568 353354 197577
rect 353298 197503 353354 197512
rect 229836 197328 229888 197334
rect 229836 197270 229888 197276
rect 229848 197033 229876 197270
rect 229834 197024 229890 197033
rect 229834 196959 229890 196968
rect 353300 194540 353352 194546
rect 353300 194482 353352 194488
rect 353312 194041 353340 194482
rect 353298 194032 353354 194041
rect 353298 193967 353354 193976
rect 230386 193216 230442 193225
rect 230386 193151 230388 193160
rect 230440 193151 230442 193160
rect 230388 193122 230440 193128
rect 230388 190460 230440 190466
rect 230388 190402 230440 190408
rect 230400 189417 230428 190402
rect 230386 189408 230442 189417
rect 230386 189343 230442 189352
rect 353300 187672 353352 187678
rect 353300 187614 353352 187620
rect 353312 186969 353340 187614
rect 353298 186960 353354 186969
rect 353298 186895 353354 186904
rect 230388 186312 230440 186318
rect 230388 186254 230440 186260
rect 230400 185609 230428 186254
rect 230386 185600 230442 185609
rect 230386 185535 230442 185544
rect 353300 183524 353352 183530
rect 353300 183466 353352 183472
rect 353312 183433 353340 183466
rect 353298 183424 353354 183433
rect 353298 183359 353354 183368
rect 229836 182164 229888 182170
rect 229836 182106 229888 182112
rect 229848 181801 229876 182106
rect 229834 181792 229890 181801
rect 229834 181727 229890 181736
rect 353300 180804 353352 180810
rect 353300 180746 353352 180752
rect 353312 179897 353340 180746
rect 353298 179888 353354 179897
rect 353298 179823 353354 179832
rect 224224 178016 224276 178022
rect 230388 178016 230440 178022
rect 224224 177958 224276 177964
rect 230386 177984 230388 177993
rect 230440 177984 230442 177993
rect 230386 177919 230442 177928
rect 353300 176656 353352 176662
rect 353300 176598 353352 176604
rect 353312 176361 353340 176598
rect 353298 176352 353354 176361
rect 353298 176287 353354 176296
rect 28264 175228 28316 175234
rect 28264 175170 28316 175176
rect 230388 175228 230440 175234
rect 230388 175170 230440 175176
rect 230400 174185 230428 175170
rect 230386 174176 230442 174185
rect 230386 174111 230442 174120
rect 353300 173868 353352 173874
rect 353300 173810 353352 173816
rect 353312 172825 353340 173810
rect 353298 172816 353354 172825
rect 353298 172751 353354 172760
rect 21364 171080 21416 171086
rect 21364 171022 21416 171028
rect 230388 171080 230440 171086
rect 230388 171022 230440 171028
rect 230400 170377 230428 171022
rect 230386 170368 230442 170377
rect 230386 170303 230442 170312
rect 13084 167000 13136 167006
rect 13084 166942 13136 166948
rect 230388 167000 230440 167006
rect 230388 166942 230440 166948
rect 353300 167000 353352 167006
rect 353300 166942 353352 166948
rect 230400 166569 230428 166942
rect 230386 166560 230442 166569
rect 230386 166495 230442 166504
rect 353312 165753 353340 166942
rect 353298 165744 353354 165753
rect 353298 165679 353354 165688
rect 3790 164656 3846 164665
rect 3790 164591 3846 164600
rect 3700 147620 3752 147626
rect 3700 147562 3752 147568
rect 3804 144906 3832 164591
rect 230388 162852 230440 162858
rect 230388 162794 230440 162800
rect 353300 162852 353352 162858
rect 353300 162794 353352 162800
rect 230400 162761 230428 162794
rect 230386 162752 230442 162761
rect 230386 162687 230442 162696
rect 353312 162217 353340 162794
rect 353298 162208 353354 162217
rect 353298 162143 353354 162152
rect 230388 160064 230440 160070
rect 230388 160006 230440 160012
rect 230400 158953 230428 160006
rect 230386 158944 230442 158953
rect 230386 158879 230442 158888
rect 353956 158681 353984 219438
rect 354048 190505 354076 364346
rect 354128 259480 354180 259486
rect 354128 259422 354180 259428
rect 354034 190496 354090 190505
rect 354034 190431 354090 190440
rect 354036 179444 354088 179450
rect 354036 179386 354088 179392
rect 353942 158672 353998 158681
rect 353942 158607 353998 158616
rect 229284 155916 229336 155922
rect 229284 155858 229336 155864
rect 353300 155916 353352 155922
rect 353300 155858 353352 155864
rect 229296 155145 229324 155858
rect 353312 155145 353340 155858
rect 229282 155136 229338 155145
rect 229282 155071 229338 155080
rect 353298 155136 353354 155145
rect 353298 155071 353354 155080
rect 353944 153264 353996 153270
rect 353944 153206 353996 153212
rect 230388 151768 230440 151774
rect 230388 151710 230440 151716
rect 353300 151768 353352 151774
rect 353300 151710 353352 151716
rect 230400 151337 230428 151710
rect 353312 151609 353340 151710
rect 353298 151600 353354 151609
rect 353298 151535 353354 151544
rect 230386 151328 230442 151337
rect 230386 151263 230442 151272
rect 230388 147620 230440 147626
rect 230388 147562 230440 147568
rect 230400 147529 230428 147562
rect 230386 147520 230442 147529
rect 230386 147455 230442 147464
rect 3792 144900 3844 144906
rect 3792 144842 3844 144848
rect 230020 144900 230072 144906
rect 230020 144842 230072 144848
rect 353300 144900 353352 144906
rect 353300 144842 353352 144848
rect 230032 143721 230060 144842
rect 353312 144537 353340 144842
rect 353298 144528 353354 144537
rect 353298 144463 353354 144472
rect 230018 143712 230074 143721
rect 230018 143647 230074 143656
rect 353956 141001 353984 153206
rect 354048 148073 354076 179386
rect 354140 169289 354168 259422
rect 355336 208214 355364 456758
rect 356716 219434 356744 509254
rect 359476 230450 359504 561682
rect 360856 251190 360884 667898
rect 579894 642152 579950 642161
rect 579894 642087 579950 642096
rect 579908 641782 579936 642087
rect 367744 641776 367796 641782
rect 367744 641718 367796 641724
rect 579896 641776 579948 641782
rect 579896 641718 579948 641724
rect 364984 535492 365036 535498
rect 364984 535434 365036 535440
rect 363604 404388 363656 404394
rect 363604 404330 363656 404336
rect 360844 251184 360896 251190
rect 360844 251126 360896 251132
rect 359464 230444 359516 230450
rect 359464 230386 359516 230392
rect 356704 219428 356756 219434
rect 356704 219370 356756 219376
rect 355324 208208 355376 208214
rect 355324 208150 355376 208156
rect 363616 198694 363644 404330
rect 364996 226302 365024 535434
rect 367756 248402 367784 641718
rect 579894 628960 579950 628969
rect 579894 628895 579950 628904
rect 579908 627978 579936 628895
rect 377404 627972 377456 627978
rect 377404 627914 377456 627920
rect 579896 627972 579948 627978
rect 579896 627914 579948 627920
rect 374644 523048 374696 523054
rect 374644 522990 374696 522996
rect 373264 430636 373316 430642
rect 373264 430578 373316 430584
rect 371884 324352 371936 324358
rect 371884 324294 371936 324300
rect 369124 271924 369176 271930
rect 369124 271866 369176 271872
rect 367744 248396 367796 248402
rect 367744 248338 367796 248344
rect 364984 226296 365036 226302
rect 364984 226238 365036 226244
rect 363604 198688 363656 198694
rect 363604 198630 363656 198636
rect 369136 173874 369164 271866
rect 371896 183530 371924 324294
rect 373276 205630 373304 430578
rect 374656 223582 374684 522990
rect 377416 244254 377444 627914
rect 580170 615768 580226 615777
rect 580170 615703 580226 615712
rect 580184 615534 580212 615703
rect 509884 615528 509936 615534
rect 509884 615470 509936 615476
rect 580172 615528 580224 615534
rect 580172 615470 580224 615476
rect 381544 416832 381596 416838
rect 381544 416774 381596 416780
rect 378784 311908 378836 311914
rect 378784 311850 378836 311856
rect 377404 244248 377456 244254
rect 377404 244190 377456 244196
rect 374644 223576 374696 223582
rect 374644 223518 374696 223524
rect 373264 205624 373316 205630
rect 373264 205566 373316 205572
rect 371884 183524 371936 183530
rect 371884 183466 371936 183472
rect 378796 180810 378824 311850
rect 381556 201482 381584 416774
rect 509896 240106 509924 615470
rect 580170 563000 580226 563009
rect 580170 562935 580226 562944
rect 580184 561746 580212 562935
rect 580172 561740 580224 561746
rect 580172 561682 580224 561688
rect 580170 536616 580226 536625
rect 580170 536551 580226 536560
rect 580184 535498 580212 536551
rect 580172 535492 580224 535498
rect 580172 535434 580224 535440
rect 580170 523424 580226 523433
rect 580170 523359 580226 523368
rect 580184 523054 580212 523359
rect 580172 523048 580224 523054
rect 580172 522990 580224 522996
rect 579618 510232 579674 510241
rect 579618 510167 579674 510176
rect 579632 509318 579660 510167
rect 579620 509312 579672 509318
rect 579620 509254 579672 509260
rect 580170 457464 580226 457473
rect 580170 457399 580226 457408
rect 580184 456822 580212 457399
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579802 431080 579858 431089
rect 579802 431015 579858 431024
rect 579816 430642 579844 431015
rect 579804 430636 579856 430642
rect 579804 430578 579856 430584
rect 579618 417888 579674 417897
rect 579618 417823 579674 417832
rect 579632 416838 579660 417823
rect 579620 416832 579672 416838
rect 579620 416774 579672 416780
rect 580170 404696 580226 404705
rect 580170 404631 580226 404640
rect 580184 404394 580212 404631
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580170 325544 580226 325553
rect 580170 325479 580226 325488
rect 580184 324358 580212 325479
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312352 580226 312361
rect 580170 312287 580226 312296
rect 580184 311914 580212 312287
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 579986 272776 580042 272785
rect 579986 272711 580042 272720
rect 580000 271930 580028 272711
rect 579988 271924 580040 271930
rect 579988 271866 580040 271872
rect 580170 259584 580226 259593
rect 580170 259519 580226 259528
rect 580184 259486 580212 259519
rect 580172 259480 580224 259486
rect 580172 259422 580224 259428
rect 580276 258074 580304 694855
rect 580354 589384 580410 589393
rect 580354 589319 580410 589328
rect 580184 258058 580304 258074
rect 580172 258052 580304 258058
rect 580224 258046 580304 258052
rect 580172 257994 580224 258000
rect 580262 246392 580318 246401
rect 580262 246327 580318 246336
rect 509884 240100 509936 240106
rect 509884 240042 509936 240048
rect 580170 220008 580226 220017
rect 580170 219943 580226 219952
rect 580184 219502 580212 219943
rect 580172 219496 580224 219502
rect 580172 219438 580224 219444
rect 381544 201476 381596 201482
rect 381544 201418 381596 201424
rect 378784 180804 378836 180810
rect 378784 180746 378836 180752
rect 579618 180432 579674 180441
rect 579618 180367 579674 180376
rect 579632 179450 579660 180367
rect 579620 179444 579672 179450
rect 579620 179386 579672 179392
rect 369124 173868 369176 173874
rect 369124 173810 369176 173816
rect 354126 169280 354182 169289
rect 354126 169215 354182 169224
rect 580276 167006 580304 246327
rect 580368 237386 580396 589319
rect 580446 576192 580502 576201
rect 580446 576127 580502 576136
rect 580356 237380 580408 237386
rect 580356 237322 580408 237328
rect 580460 233238 580488 576127
rect 580538 483848 580594 483857
rect 580538 483783 580594 483792
rect 580448 233232 580500 233238
rect 580354 233200 580410 233209
rect 580448 233174 580500 233180
rect 580354 233135 580410 233144
rect 580264 167000 580316 167006
rect 580264 166942 580316 166948
rect 580368 162858 580396 233135
rect 580552 215286 580580 483783
rect 580630 470656 580686 470665
rect 580630 470591 580686 470600
rect 580540 215280 580592 215286
rect 580540 215222 580592 215228
rect 580644 212498 580672 470591
rect 580722 378312 580778 378321
rect 580722 378247 580778 378256
rect 580632 212492 580684 212498
rect 580632 212434 580684 212440
rect 580446 206816 580502 206825
rect 580446 206751 580502 206760
rect 580356 162852 580408 162858
rect 580356 162794 580408 162800
rect 580460 155922 580488 206751
rect 580736 194546 580764 378247
rect 580814 351928 580870 351937
rect 580814 351863 580870 351872
rect 580724 194540 580776 194546
rect 580724 194482 580776 194488
rect 580538 193624 580594 193633
rect 580538 193559 580594 193568
rect 580448 155916 580500 155922
rect 580448 155858 580500 155864
rect 579618 154048 579674 154057
rect 579618 153983 579674 153992
rect 579632 153270 579660 153983
rect 579620 153264 579672 153270
rect 579620 153206 579672 153212
rect 580552 151774 580580 193559
rect 580828 187678 580856 351863
rect 580906 299160 580962 299169
rect 580906 299095 580962 299104
rect 580816 187672 580868 187678
rect 580816 187614 580868 187620
rect 580920 176662 580948 299095
rect 580908 176656 580960 176662
rect 580908 176598 580960 176604
rect 580630 167240 580686 167249
rect 580630 167175 580686 167184
rect 580540 151768 580592 151774
rect 580540 151710 580592 151716
rect 354034 148064 354090 148073
rect 354034 147999 354090 148008
rect 580644 144906 580672 167175
rect 580632 144900 580684 144906
rect 580632 144842 580684 144848
rect 353942 140992 353998 141001
rect 353942 140927 353998 140936
rect 580170 140856 580226 140865
rect 353300 140820 353352 140826
rect 580170 140791 580172 140800
rect 353300 140762 353352 140768
rect 580224 140791 580226 140800
rect 580172 140762 580224 140768
rect 3424 140752 3476 140758
rect 3424 140694 3476 140700
rect 230388 140752 230440 140758
rect 230388 140694 230440 140700
rect 230400 139913 230428 140694
rect 230386 139904 230442 139913
rect 230386 139839 230442 139848
rect 3422 138816 3478 138825
rect 3422 138751 3478 138760
rect 3436 136610 3464 138751
rect 353312 137465 353340 140762
rect 353298 137456 353354 137465
rect 353298 137391 353354 137400
rect 3424 136604 3476 136610
rect 3424 136546 3476 136552
rect 229652 136604 229704 136610
rect 229652 136546 229704 136552
rect 229664 136105 229692 136546
rect 229650 136096 229706 136105
rect 229650 136031 229706 136040
rect 354218 133920 354274 133929
rect 354218 133855 354274 133864
rect 229742 132288 229798 132297
rect 229742 132223 229798 132232
rect 3608 128376 3660 128382
rect 3608 128318 3660 128324
rect 3516 116000 3568 116006
rect 3516 115942 3568 115948
rect 3148 113144 3200 113150
rect 3148 113086 3200 113092
rect 3160 112985 3188 113086
rect 3146 112976 3202 112985
rect 3146 112911 3202 112920
rect 3424 104916 3476 104922
rect 3424 104858 3476 104864
rect 3332 88324 3384 88330
rect 3332 88266 3384 88272
rect 3344 87145 3372 88266
rect 3330 87136 3386 87145
rect 3330 87071 3386 87080
rect 3332 74520 3384 74526
rect 3332 74462 3384 74468
rect 3344 74225 3372 74462
rect 3330 74216 3386 74225
rect 3330 74151 3386 74160
rect 3240 49700 3292 49706
rect 3240 49642 3292 49648
rect 3252 48385 3280 49642
rect 3238 48376 3294 48385
rect 3238 48311 3294 48320
rect 3332 35896 3384 35902
rect 3332 35838 3384 35844
rect 3344 35465 3372 35838
rect 3330 35456 3386 35465
rect 3330 35391 3386 35400
rect 3436 22545 3464 104858
rect 3528 61305 3556 115942
rect 3620 100065 3648 128318
rect 229756 113150 229784 132223
rect 353942 130384 353998 130393
rect 353942 130319 353998 130328
rect 230386 128480 230442 128489
rect 230386 128415 230442 128424
rect 230400 128382 230428 128415
rect 230388 128376 230440 128382
rect 230388 128318 230440 128324
rect 230110 124672 230166 124681
rect 230110 124607 230166 124616
rect 230018 120864 230074 120873
rect 230018 120799 230074 120808
rect 229926 113248 229982 113257
rect 229926 113183 229982 113192
rect 229744 113144 229796 113150
rect 229744 113086 229796 113092
rect 229834 109440 229890 109449
rect 229834 109375 229890 109384
rect 229742 101824 229798 101833
rect 229742 101759 229798 101768
rect 3606 100056 3662 100065
rect 3606 99991 3662 100000
rect 128360 97504 128412 97510
rect 128360 97446 128412 97452
rect 121460 97368 121512 97374
rect 121460 97310 121512 97316
rect 28264 97300 28316 97306
rect 28264 97242 28316 97248
rect 26240 75200 26292 75206
rect 26240 75142 26292 75148
rect 20720 66904 20772 66910
rect 20720 66846 20772 66852
rect 3514 61296 3570 61305
rect 3514 61231 3570 61240
rect 3422 22536 3478 22545
rect 3422 22471 3478 22480
rect 3424 9648 3476 9654
rect 3422 9616 3424 9625
rect 3476 9616 3478 9625
rect 3422 9551 3478 9560
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 19812 480 19840 6122
rect 20732 2378 20760 66846
rect 22100 54528 22152 54534
rect 22100 54470 22152 54476
rect 22112 16574 22140 54470
rect 26252 16574 26280 75142
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 27632 16574 27660 21354
rect 22112 16546 23152 16574
rect 26252 16546 26464 16574
rect 27632 16546 28212 16574
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20916 480 20944 6190
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 22020 480 22048 2314
rect 23124 480 23152 16546
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 24214 3360 24270 3369
rect 24214 3295 24270 3304
rect 24228 480 24256 3295
rect 25332 480 25360 3878
rect 26436 480 26464 16546
rect 28184 3482 28212 16546
rect 28276 3942 28304 97242
rect 81440 96008 81492 96014
rect 81440 95950 81492 95956
rect 75920 95940 75972 95946
rect 75920 95882 75972 95888
rect 66260 94580 66312 94586
rect 66260 94522 66312 94528
rect 40040 94512 40092 94518
rect 40040 94454 40092 94460
rect 30380 84856 30432 84862
rect 30380 84798 30432 84804
rect 30392 16574 30420 84798
rect 35900 76560 35952 76566
rect 35900 76502 35952 76508
rect 35164 61396 35216 61402
rect 35164 61338 35216 61344
rect 31760 46232 31812 46238
rect 31760 46174 31812 46180
rect 31772 16574 31800 46174
rect 34520 32428 34572 32434
rect 34520 32370 34572 32376
rect 32404 31068 32456 31074
rect 32404 31010 32456 31016
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 28264 3936 28316 3942
rect 28264 3878 28316 3884
rect 28184 3454 28672 3482
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 27540 480 27568 2994
rect 28644 480 28672 3454
rect 29736 3460 29788 3466
rect 29736 3402 29788 3408
rect 29748 480 29776 3402
rect 30852 480 30880 16546
rect 31956 480 31984 16546
rect 32416 3058 32444 31010
rect 34532 16574 34560 32370
rect 34532 16546 35112 16574
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 33060 480 33088 3538
rect 34152 3528 34204 3534
rect 34152 3470 34204 3476
rect 35084 3482 35112 16546
rect 35176 3602 35204 61338
rect 35912 16574 35940 76502
rect 38660 37936 38712 37942
rect 38660 37878 38712 37884
rect 38672 16574 38700 37878
rect 40052 16574 40080 94454
rect 63500 93220 63552 93226
rect 63500 93162 63552 93168
rect 56600 93152 56652 93158
rect 56600 93094 56652 93100
rect 53840 83496 53892 83502
rect 53840 83438 53892 83444
rect 42800 82136 42852 82142
rect 42800 82078 42852 82084
rect 35912 16546 36400 16574
rect 38672 16546 39712 16574
rect 40052 16546 40816 16574
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 34164 480 34192 3470
rect 35084 3454 35296 3482
rect 35268 480 35296 3454
rect 36372 480 36400 16546
rect 38568 3664 38620 3670
rect 38568 3606 38620 3612
rect 37464 3392 37516 3398
rect 37464 3334 37516 3340
rect 37476 480 37504 3334
rect 38580 480 38608 3606
rect 39684 480 39712 16546
rect 40788 480 40816 16546
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 41892 480 41920 3674
rect 42812 3602 42840 82078
rect 46940 72480 46992 72486
rect 46940 72422 46992 72428
rect 44180 36576 44232 36582
rect 44180 36518 44232 36524
rect 44192 16574 44220 36518
rect 46952 16574 46980 72422
rect 49700 64184 49752 64190
rect 49700 64126 49752 64132
rect 48320 33788 48372 33794
rect 48320 33730 48372 33736
rect 48332 16574 48360 33730
rect 49712 16574 49740 64126
rect 44192 16546 45232 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50752 16574
rect 42984 3800 43036 3806
rect 42984 3742 43036 3748
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 42996 480 43024 3742
rect 44272 3664 44324 3670
rect 44272 3606 44324 3612
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 44100 480 44128 3538
rect 44284 3398 44312 3606
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 45204 480 45232 16546
rect 46296 3868 46348 3874
rect 46296 3810 46348 3816
rect 46308 480 46336 3810
rect 47412 480 47440 16546
rect 48516 480 48544 16546
rect 49608 3936 49660 3942
rect 49608 3878 49660 3884
rect 49620 480 49648 3878
rect 50724 480 50752 16546
rect 51816 10328 51868 10334
rect 51816 10270 51868 10276
rect 51828 480 51856 10270
rect 52920 4004 52972 4010
rect 52920 3946 52972 3952
rect 52932 480 52960 3946
rect 53852 3398 53880 83438
rect 53932 55888 53984 55894
rect 53932 55830 53984 55836
rect 53944 16574 53972 55830
rect 56612 16574 56640 93094
rect 57980 68332 58032 68338
rect 57980 68274 58032 68280
rect 57992 16574 58020 68274
rect 59360 65544 59412 65550
rect 59360 65486 59412 65492
rect 53944 16546 54064 16574
rect 56612 16546 57376 16574
rect 57992 16546 58480 16574
rect 53840 3392 53892 3398
rect 53840 3334 53892 3340
rect 54036 480 54064 16546
rect 56232 4072 56284 4078
rect 56232 4014 56284 4020
rect 55128 3392 55180 3398
rect 55128 3334 55180 3340
rect 55140 480 55168 3334
rect 56244 480 56272 4014
rect 57348 480 57376 16546
rect 58452 480 58480 16546
rect 59372 3398 59400 65486
rect 60740 22772 60792 22778
rect 60740 22714 60792 22720
rect 60752 16574 60780 22714
rect 63512 16574 63540 93162
rect 64880 29640 64932 29646
rect 64880 29582 64932 29588
rect 64892 16574 64920 29582
rect 66272 16574 66300 94522
rect 70400 83564 70452 83570
rect 70400 83506 70452 83512
rect 67640 51740 67692 51746
rect 67640 51682 67692 51688
rect 67652 16574 67680 51682
rect 60752 16546 61792 16574
rect 63512 16546 64000 16574
rect 64892 16546 65104 16574
rect 66272 16546 67312 16574
rect 67652 16546 68416 16574
rect 59544 4140 59596 4146
rect 59544 4082 59596 4088
rect 59360 3392 59412 3398
rect 59360 3334 59412 3340
rect 59556 480 59584 4082
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60660 480 60688 3334
rect 61764 480 61792 16546
rect 62856 3392 62908 3398
rect 62856 3334 62908 3340
rect 62868 480 62896 3334
rect 63972 480 64000 16546
rect 65076 480 65104 16546
rect 66168 7608 66220 7614
rect 66168 7550 66220 7556
rect 66180 480 66208 7550
rect 67284 480 67312 16546
rect 68388 480 68416 16546
rect 69480 11756 69532 11762
rect 69480 11698 69532 11704
rect 69492 480 69520 11698
rect 70412 3482 70440 83506
rect 70492 53100 70544 53106
rect 70492 53042 70544 53048
rect 70504 4214 70532 53042
rect 74540 50380 74592 50386
rect 74540 50322 74592 50328
rect 71780 19984 71832 19990
rect 71780 19926 71832 19932
rect 71792 16574 71820 19926
rect 73160 17264 73212 17270
rect 73160 17206 73212 17212
rect 73172 16574 73200 17206
rect 74552 16574 74580 50322
rect 71792 16546 72832 16574
rect 73172 16546 73936 16574
rect 74552 16546 75040 16574
rect 70492 4208 70544 4214
rect 70492 4150 70544 4156
rect 71688 4208 71740 4214
rect 71688 4150 71740 4156
rect 70412 3454 70624 3482
rect 70596 480 70624 3454
rect 71700 480 71728 4150
rect 72804 480 72832 16546
rect 73908 480 73936 16546
rect 75012 480 75040 16546
rect 75932 3330 75960 95882
rect 80060 89004 80112 89010
rect 80060 88946 80112 88952
rect 78680 77988 78732 77994
rect 78680 77930 78732 77936
rect 77300 28280 77352 28286
rect 77300 28222 77352 28228
rect 76012 18624 76064 18630
rect 76012 18566 76064 18572
rect 76024 16574 76052 18566
rect 77312 16574 77340 28222
rect 78692 16574 78720 77930
rect 80072 16574 80100 88946
rect 76024 16546 76144 16574
rect 77312 16546 78352 16574
rect 78692 16546 79456 16574
rect 80072 16546 80560 16574
rect 75920 3324 75972 3330
rect 75920 3266 75972 3272
rect 76116 480 76144 16546
rect 77208 3324 77260 3330
rect 77208 3266 77260 3272
rect 77220 480 77248 3266
rect 78324 480 78352 16546
rect 79428 480 79456 16546
rect 80532 480 80560 16546
rect 81452 3330 81480 95950
rect 106280 91792 106332 91798
rect 106280 91734 106332 91740
rect 92480 90364 92532 90370
rect 92480 90306 92532 90312
rect 89720 86284 89772 86290
rect 89720 86226 89772 86232
rect 88340 84924 88392 84930
rect 88340 84866 88392 84872
rect 82820 76628 82872 76634
rect 82820 76570 82872 76576
rect 81532 26920 81584 26926
rect 81532 26862 81584 26868
rect 81544 16574 81572 26862
rect 82832 16574 82860 76570
rect 86960 68400 87012 68406
rect 86960 68342 87012 68348
rect 84200 39364 84252 39370
rect 84200 39306 84252 39312
rect 84212 16574 84240 39306
rect 81544 16546 81664 16574
rect 82832 16546 83872 16574
rect 84212 16546 84976 16574
rect 81440 3324 81492 3330
rect 81440 3266 81492 3272
rect 81636 480 81664 16546
rect 82728 3324 82780 3330
rect 82728 3266 82780 3272
rect 82740 480 82768 3266
rect 83844 480 83872 16546
rect 84948 480 84976 16546
rect 86040 4820 86092 4826
rect 86040 4762 86092 4768
rect 86052 480 86080 4762
rect 86972 3482 87000 68342
rect 87052 24132 87104 24138
rect 87052 24074 87104 24080
rect 87064 4214 87092 24074
rect 88352 16574 88380 84866
rect 89732 16574 89760 86226
rect 91100 73840 91152 73846
rect 91100 73782 91152 73788
rect 91112 16574 91140 73782
rect 88352 16546 89392 16574
rect 89732 16546 90496 16574
rect 91112 16546 91600 16574
rect 87052 4208 87104 4214
rect 87052 4150 87104 4156
rect 88248 4208 88300 4214
rect 88248 4150 88300 4156
rect 86972 3454 87184 3482
rect 87156 480 87184 3454
rect 88260 480 88288 4150
rect 89364 480 89392 16546
rect 90468 480 90496 16546
rect 91572 480 91600 16546
rect 92492 3330 92520 90306
rect 98000 89072 98052 89078
rect 98000 89014 98052 89020
rect 96620 79348 96672 79354
rect 96620 79290 96672 79296
rect 93860 47592 93912 47598
rect 93860 47534 93912 47540
rect 92572 32496 92624 32502
rect 92572 32438 92624 32444
rect 92584 16574 92612 32438
rect 93872 16574 93900 47534
rect 95240 31136 95292 31142
rect 95240 31078 95292 31084
rect 95252 16574 95280 31078
rect 96632 16574 96660 79290
rect 92584 16546 92704 16574
rect 93872 16546 94912 16574
rect 95252 16546 96016 16574
rect 96632 16546 97120 16574
rect 92480 3324 92532 3330
rect 92480 3266 92532 3272
rect 92676 480 92704 16546
rect 93768 3324 93820 3330
rect 93768 3266 93820 3272
rect 93780 480 93808 3266
rect 94884 480 94912 16546
rect 95988 480 96016 16546
rect 97092 480 97120 16546
rect 98012 3330 98040 89014
rect 99380 78056 99432 78062
rect 99380 77998 99432 78004
rect 98092 25560 98144 25566
rect 98092 25502 98144 25508
rect 98104 16574 98132 25502
rect 99392 16574 99420 77998
rect 103520 75268 103572 75274
rect 103520 75210 103572 75216
rect 102140 29708 102192 29714
rect 102140 29650 102192 29656
rect 102152 16574 102180 29650
rect 98104 16546 98224 16574
rect 99392 16546 100432 16574
rect 102152 16546 102640 16574
rect 98000 3324 98052 3330
rect 98000 3266 98052 3272
rect 98196 480 98224 16546
rect 99288 3324 99340 3330
rect 99288 3266 99340 3272
rect 99300 480 99328 3266
rect 100404 480 100432 16546
rect 101496 15904 101548 15910
rect 101496 15846 101548 15852
rect 101508 480 101536 15846
rect 102612 480 102640 16546
rect 103532 3330 103560 75210
rect 103612 62824 103664 62830
rect 103612 62766 103664 62772
rect 103624 16574 103652 62766
rect 106292 16574 106320 91734
rect 115940 87644 115992 87650
rect 115940 87586 115992 87592
rect 109040 71052 109092 71058
rect 109040 70994 109092 71000
rect 107660 44872 107712 44878
rect 107660 44814 107712 44820
rect 107672 16574 107700 44814
rect 103624 16546 103744 16574
rect 106292 16546 107056 16574
rect 107672 16546 108160 16574
rect 103520 3324 103572 3330
rect 103520 3266 103572 3272
rect 103716 480 103744 16546
rect 105912 9172 105964 9178
rect 105912 9114 105964 9120
rect 104808 3324 104860 3330
rect 104808 3266 104860 3272
rect 104820 480 104848 3266
rect 105924 480 105952 9114
rect 107028 480 107056 16546
rect 108132 480 108160 16546
rect 109052 3330 109080 70994
rect 113180 69692 113232 69698
rect 113180 69634 113232 69640
rect 110420 40724 110472 40730
rect 110420 40666 110472 40672
rect 109132 17332 109184 17338
rect 109132 17274 109184 17280
rect 109144 16574 109172 17274
rect 110432 16574 110460 40666
rect 111800 28348 111852 28354
rect 111800 28290 111852 28296
rect 111812 16574 111840 28290
rect 113192 16574 113220 69634
rect 114560 66972 114612 66978
rect 114560 66914 114612 66920
rect 109144 16546 109264 16574
rect 110432 16546 111472 16574
rect 111812 16546 112576 16574
rect 113192 16546 113680 16574
rect 109040 3324 109092 3330
rect 109040 3266 109092 3272
rect 109236 480 109264 16546
rect 110328 3324 110380 3330
rect 110328 3266 110380 3272
rect 110340 480 110368 3266
rect 111444 480 111472 16546
rect 112548 480 112576 16546
rect 113652 480 113680 16546
rect 114572 3482 114600 66914
rect 114652 26988 114704 26994
rect 114652 26930 114704 26936
rect 114664 4214 114692 26930
rect 115952 16574 115980 87586
rect 120080 80708 120132 80714
rect 120080 80650 120132 80656
rect 117320 42084 117372 42090
rect 117320 42026 117372 42032
rect 117332 16574 117360 42026
rect 118700 24200 118752 24206
rect 118700 24142 118752 24148
rect 118712 16574 118740 24142
rect 115952 16546 116992 16574
rect 117332 16546 118096 16574
rect 118712 16546 119200 16574
rect 114652 4208 114704 4214
rect 114652 4150 114704 4156
rect 115848 4208 115900 4214
rect 115848 4150 115900 4156
rect 114572 3454 114784 3482
rect 114756 480 114784 3454
rect 115860 480 115888 4150
rect 116964 480 116992 16546
rect 118068 480 118096 16546
rect 119172 480 119200 16546
rect 120092 3482 120120 80650
rect 120172 43444 120224 43450
rect 120172 43386 120224 43392
rect 120184 4214 120212 43386
rect 121472 16574 121500 97310
rect 122840 61464 122892 61470
rect 122840 61406 122892 61412
rect 122852 16574 122880 61406
rect 125600 60036 125652 60042
rect 125600 59978 125652 59984
rect 121472 16546 122512 16574
rect 122852 16546 123616 16574
rect 120172 4208 120224 4214
rect 120172 4150 120224 4156
rect 121368 4208 121420 4214
rect 121368 4150 121420 4156
rect 120092 3454 120304 3482
rect 120276 480 120304 3454
rect 121380 480 121408 4150
rect 122484 480 122512 16546
rect 123588 480 123616 16546
rect 124680 14476 124732 14482
rect 124680 14418 124732 14424
rect 124692 480 124720 14418
rect 125612 3330 125640 59978
rect 125692 25628 125744 25634
rect 125692 25570 125744 25576
rect 125704 16574 125732 25570
rect 128372 16574 128400 97446
rect 224960 96280 225012 96286
rect 224960 96222 225012 96228
rect 216680 96212 216732 96218
rect 216680 96154 216732 96160
rect 195980 96144 196032 96150
rect 195980 96086 196032 96092
rect 169760 96076 169812 96082
rect 169760 96018 169812 96024
rect 155960 91860 156012 91866
rect 155960 91802 156012 91808
rect 136640 89140 136692 89146
rect 136640 89082 136692 89088
rect 129740 58676 129792 58682
rect 129740 58618 129792 58624
rect 129752 16574 129780 58618
rect 132500 57248 132552 57254
rect 132500 57190 132552 57196
rect 131120 49020 131172 49026
rect 131120 48962 131172 48968
rect 131132 16574 131160 48962
rect 132512 16574 132540 57190
rect 133880 35216 133932 35222
rect 133880 35158 133932 35164
rect 133892 16574 133920 35158
rect 125704 16546 125824 16574
rect 128372 16546 129136 16574
rect 129752 16546 130240 16574
rect 131132 16546 131344 16574
rect 132512 16546 133552 16574
rect 133892 16546 134656 16574
rect 125600 3324 125652 3330
rect 125600 3266 125652 3272
rect 125796 480 125824 16546
rect 127992 13116 128044 13122
rect 127992 13058 128044 13064
rect 126888 3324 126940 3330
rect 126888 3266 126940 3272
rect 126900 480 126928 3266
rect 128004 480 128032 13058
rect 129108 480 129136 16546
rect 130212 480 130240 16546
rect 131316 480 131344 16546
rect 132408 3324 132460 3330
rect 132408 3266 132460 3272
rect 132420 480 132448 3266
rect 133524 480 133552 16546
rect 134628 480 134656 16546
rect 135720 3256 135772 3262
rect 135720 3198 135772 3204
rect 135732 480 135760 3198
rect 136652 2786 136680 89082
rect 139400 86352 139452 86358
rect 139400 86294 139452 86300
rect 138020 82204 138072 82210
rect 138020 82146 138072 82152
rect 138032 16574 138060 82146
rect 139412 16574 139440 86294
rect 149060 84992 149112 84998
rect 149060 84934 149112 84940
rect 142160 80776 142212 80782
rect 142160 80718 142212 80724
rect 140780 65612 140832 65618
rect 140780 65554 140832 65560
rect 140792 16574 140820 65554
rect 138032 16546 139072 16574
rect 139412 16546 140176 16574
rect 140792 16546 141280 16574
rect 136824 4956 136876 4962
rect 136824 4898 136876 4904
rect 136640 2780 136692 2786
rect 136640 2722 136692 2728
rect 136836 480 136864 4898
rect 137928 2780 137980 2786
rect 137928 2722 137980 2728
rect 137940 480 137968 2722
rect 139044 480 139072 16546
rect 140148 480 140176 16546
rect 141252 480 141280 16546
rect 142172 3194 142200 80718
rect 146300 79416 146352 79422
rect 146300 79358 146352 79364
rect 143540 62892 143592 62898
rect 143540 62834 143592 62840
rect 142252 43512 142304 43518
rect 142252 43454 142304 43460
rect 142264 16574 142292 43454
rect 143552 16574 143580 62834
rect 144920 36644 144972 36650
rect 144920 36586 144972 36592
rect 144932 16574 144960 36586
rect 146312 16574 146340 79358
rect 147680 60104 147732 60110
rect 147680 60046 147732 60052
rect 142264 16546 142384 16574
rect 143552 16546 144592 16574
rect 144932 16546 145696 16574
rect 146312 16546 146800 16574
rect 142160 3188 142212 3194
rect 142160 3130 142212 3136
rect 142356 480 142384 16546
rect 143448 3188 143500 3194
rect 143448 3130 143500 3136
rect 143460 480 143488 3130
rect 144564 480 144592 16546
rect 145668 480 145696 16546
rect 146772 480 146800 16546
rect 147692 3482 147720 60046
rect 147772 18692 147824 18698
rect 147772 18634 147824 18640
rect 147784 4214 147812 18634
rect 149072 16574 149100 84934
rect 153200 78124 153252 78130
rect 153200 78066 153252 78072
rect 150440 58744 150492 58750
rect 150440 58686 150492 58692
rect 150452 16574 150480 58686
rect 151820 33856 151872 33862
rect 151820 33798 151872 33804
rect 151832 16574 151860 33798
rect 149072 16546 150112 16574
rect 150452 16546 151216 16574
rect 151832 16546 152320 16574
rect 147772 4208 147824 4214
rect 147772 4150 147824 4156
rect 148968 4208 149020 4214
rect 148968 4150 149020 4156
rect 147692 3454 147904 3482
rect 147876 480 147904 3454
rect 148980 480 149008 4150
rect 150084 480 150112 16546
rect 151188 480 151216 16546
rect 152292 480 152320 16546
rect 153212 3482 153240 78066
rect 153292 72548 153344 72554
rect 153292 72490 153344 72496
rect 153304 4214 153332 72490
rect 154580 20052 154632 20058
rect 154580 19994 154632 20000
rect 154592 16574 154620 19994
rect 155972 16574 156000 91802
rect 158720 83632 158772 83638
rect 158720 83574 158772 83580
rect 157340 57316 157392 57322
rect 157340 57258 157392 57264
rect 157352 16574 157380 57258
rect 154592 16546 155632 16574
rect 155972 16546 156736 16574
rect 157352 16546 157840 16574
rect 153292 4208 153344 4214
rect 153292 4150 153344 4156
rect 154488 4208 154540 4214
rect 154488 4150 154540 4156
rect 153212 3454 153424 3482
rect 153396 480 153424 3454
rect 154500 480 154528 4150
rect 155604 480 155632 16546
rect 156708 480 156736 16546
rect 157812 480 157840 16546
rect 158732 3194 158760 83574
rect 165620 82272 165672 82278
rect 165620 82214 165672 82220
rect 162860 76696 162912 76702
rect 162860 76638 162912 76644
rect 161480 64252 161532 64258
rect 161480 64194 161532 64200
rect 160100 55956 160152 55962
rect 160100 55898 160152 55904
rect 160112 16574 160140 55898
rect 161492 16574 161520 64194
rect 162872 16574 162900 76638
rect 164240 54596 164292 54602
rect 164240 54538 164292 54544
rect 160112 16546 161152 16574
rect 161492 16546 162256 16574
rect 162872 16546 163360 16574
rect 158904 11824 158956 11830
rect 158904 11766 158956 11772
rect 158720 3188 158772 3194
rect 158720 3130 158772 3136
rect 158916 480 158944 11766
rect 160008 3188 160060 3194
rect 160008 3130 160060 3136
rect 160020 480 160048 3130
rect 161124 480 161152 16546
rect 162228 480 162256 16546
rect 163332 480 163360 16546
rect 164252 3482 164280 54538
rect 164332 21480 164384 21486
rect 164332 21422 164384 21428
rect 164344 4214 164372 21422
rect 165632 16574 165660 82214
rect 167000 53168 167052 53174
rect 167000 53110 167052 53116
rect 167012 16574 167040 53110
rect 168380 22840 168432 22846
rect 168380 22782 168432 22788
rect 168392 16574 168420 22782
rect 165632 16546 166672 16574
rect 167012 16546 167776 16574
rect 168392 16546 168880 16574
rect 164332 4208 164384 4214
rect 164332 4150 164384 4156
rect 165528 4208 165580 4214
rect 165528 4150 165580 4156
rect 164252 3454 164464 3482
rect 164436 480 164464 3454
rect 165540 480 165568 4150
rect 166644 480 166672 16546
rect 167748 480 167776 16546
rect 168852 480 168880 16546
rect 169772 3482 169800 96018
rect 175280 94648 175332 94654
rect 175280 94590 175332 94596
rect 173900 90432 173952 90438
rect 173900 90374 173952 90380
rect 169852 75336 169904 75342
rect 169852 75278 169904 75284
rect 169864 4214 169892 75278
rect 171140 61532 171192 61538
rect 171140 61474 171192 61480
rect 171152 16574 171180 61474
rect 173912 16574 173940 90374
rect 171152 16546 172192 16574
rect 173912 16546 174400 16574
rect 169852 4208 169904 4214
rect 169852 4150 169904 4156
rect 171048 4208 171100 4214
rect 171048 4150 171100 4156
rect 169772 3454 169984 3482
rect 169956 480 169984 3454
rect 171060 480 171088 4150
rect 172164 480 172192 16546
rect 173256 7676 173308 7682
rect 173256 7618 173308 7624
rect 173268 480 173296 7618
rect 174372 480 174400 16546
rect 175292 3194 175320 94590
rect 179420 93288 179472 93294
rect 179420 93230 179472 93236
rect 176660 72616 176712 72622
rect 176660 72558 176712 72564
rect 175372 51808 175424 51814
rect 175372 51750 175424 51756
rect 175384 16574 175412 51750
rect 176672 16574 176700 72558
rect 178040 50448 178092 50454
rect 178040 50390 178092 50396
rect 178052 16574 178080 50390
rect 179432 16574 179460 93230
rect 182180 91928 182232 91934
rect 182180 91870 182232 91876
rect 180800 71120 180852 71126
rect 180800 71062 180852 71068
rect 175384 16546 175504 16574
rect 176672 16546 177712 16574
rect 178052 16546 178816 16574
rect 179432 16546 179920 16574
rect 175280 3188 175332 3194
rect 175280 3130 175332 3136
rect 175476 480 175504 16546
rect 176568 3188 176620 3194
rect 176568 3130 176620 3136
rect 176580 480 176608 3130
rect 177684 480 177712 16546
rect 178788 480 178816 16546
rect 179892 480 179920 16546
rect 180812 3482 180840 71062
rect 180892 47660 180944 47666
rect 180892 47602 180944 47608
rect 180904 4214 180932 47602
rect 182192 16574 182220 91870
rect 189080 90500 189132 90506
rect 189080 90442 189132 90448
rect 187700 87712 187752 87718
rect 187700 87654 187752 87660
rect 183560 69760 183612 69766
rect 183560 69702 183612 69708
rect 183572 16574 183600 69702
rect 186320 68468 186372 68474
rect 186320 68410 186372 68416
rect 184940 46300 184992 46306
rect 184940 46242 184992 46248
rect 184952 16574 184980 46242
rect 182192 16546 183232 16574
rect 183572 16546 184336 16574
rect 184952 16546 185440 16574
rect 180892 4208 180944 4214
rect 180892 4150 180944 4156
rect 182088 4208 182140 4214
rect 182088 4150 182140 4156
rect 180812 3454 181024 3482
rect 180996 480 181024 3454
rect 182100 480 182128 4150
rect 183204 480 183232 16546
rect 184308 480 184336 16546
rect 185412 480 185440 16546
rect 186332 3194 186360 68410
rect 187712 16574 187740 87654
rect 189092 16574 189120 90442
rect 191840 89208 191892 89214
rect 191840 89150 191892 89156
rect 190460 80844 190512 80850
rect 190460 80786 190512 80792
rect 190472 16574 190500 80786
rect 187712 16546 188752 16574
rect 189092 16546 189856 16574
rect 190472 16546 190960 16574
rect 186504 10396 186556 10402
rect 186504 10338 186556 10344
rect 186320 3188 186372 3194
rect 186320 3130 186372 3136
rect 186516 480 186544 10338
rect 187608 3188 187660 3194
rect 187608 3130 187660 3136
rect 187620 480 187648 3130
rect 188724 480 188752 16546
rect 189828 480 189856 16546
rect 190932 480 190960 16546
rect 191852 3194 191880 89150
rect 193220 67040 193272 67046
rect 193220 66982 193272 66988
rect 191932 44940 191984 44946
rect 191932 44882 191984 44888
rect 191944 16574 191972 44882
rect 193232 16574 193260 66982
rect 195992 16574 196020 96086
rect 213920 94784 213972 94790
rect 213920 94726 213972 94732
rect 198740 94716 198792 94722
rect 198740 94658 198792 94664
rect 197360 86420 197412 86426
rect 197360 86362 197412 86368
rect 191944 16546 192064 16574
rect 193232 16546 194272 16574
rect 195992 16546 196480 16574
rect 191840 3188 191892 3194
rect 191840 3130 191892 3136
rect 192036 480 192064 16546
rect 193128 3188 193180 3194
rect 193128 3130 193180 3136
rect 193140 480 193168 3130
rect 194244 480 194272 16546
rect 195336 13184 195388 13190
rect 195336 13126 195388 13132
rect 195348 480 195376 13126
rect 196452 480 196480 16546
rect 197372 3482 197400 86362
rect 197452 71188 197504 71194
rect 197452 71130 197504 71136
rect 197464 4214 197492 71130
rect 198752 16574 198780 94658
rect 205640 93356 205692 93362
rect 205640 93298 205692 93304
rect 202880 85060 202932 85066
rect 202880 85002 202932 85008
rect 200120 73908 200172 73914
rect 200120 73850 200172 73856
rect 200132 16574 200160 73850
rect 201500 69828 201552 69834
rect 201500 69770 201552 69776
rect 201512 16574 201540 69770
rect 198752 16546 199792 16574
rect 200132 16546 200896 16574
rect 201512 16546 202000 16574
rect 197452 4208 197504 4214
rect 197452 4150 197504 4156
rect 198648 4208 198700 4214
rect 198648 4150 198700 4156
rect 197372 3454 197584 3482
rect 197556 480 197584 3454
rect 198660 480 198688 4150
rect 199764 480 199792 16546
rect 200868 480 200896 16546
rect 201972 480 202000 16546
rect 202892 3482 202920 85002
rect 202972 79484 203024 79490
rect 202972 79426 203024 79432
rect 202984 4214 203012 79426
rect 204260 42152 204312 42158
rect 204260 42094 204312 42100
rect 204272 16574 204300 42094
rect 205652 16574 205680 93298
rect 212540 91996 212592 92002
rect 212540 91938 212592 91944
rect 208400 87780 208452 87786
rect 208400 87722 208452 87728
rect 207020 78192 207072 78198
rect 207020 78134 207072 78140
rect 207032 16574 207060 78134
rect 204272 16546 205312 16574
rect 205652 16546 206416 16574
rect 207032 16546 207520 16574
rect 202972 4208 203024 4214
rect 202972 4150 203024 4156
rect 204168 4208 204220 4214
rect 204168 4150 204220 4156
rect 202892 3454 203104 3482
rect 203076 480 203104 3454
rect 204180 480 204208 4150
rect 205284 480 205312 16546
rect 206388 480 206416 16546
rect 207492 480 207520 16546
rect 208412 3194 208440 87722
rect 209780 64320 209832 64326
rect 209780 64262 209832 64268
rect 209792 16574 209820 64262
rect 211160 40792 211212 40798
rect 211160 40734 211212 40740
rect 211172 16574 211200 40734
rect 212552 16574 212580 91938
rect 209792 16546 210832 16574
rect 211172 16546 211936 16574
rect 212552 16546 213040 16574
rect 208584 14544 208636 14550
rect 208584 14486 208636 14492
rect 208400 3188 208452 3194
rect 208400 3130 208452 3136
rect 208596 480 208624 14486
rect 209688 3188 209740 3194
rect 209688 3130 209740 3136
rect 209700 480 209728 3130
rect 210804 480 210832 16546
rect 211908 480 211936 16546
rect 213012 480 213040 16546
rect 213932 3482 213960 94726
rect 215300 83700 215352 83706
rect 215300 83642 215352 83648
rect 214012 65680 214064 65686
rect 214012 65622 214064 65628
rect 214024 4214 214052 65622
rect 215312 16574 215340 83642
rect 216692 16574 216720 96154
rect 219440 93424 219492 93430
rect 219440 93366 219492 93372
rect 218060 39432 218112 39438
rect 218060 39374 218112 39380
rect 218072 16574 218100 39374
rect 215312 16546 216352 16574
rect 216692 16546 217456 16574
rect 218072 16546 218560 16574
rect 214012 4208 214064 4214
rect 214012 4150 214064 4156
rect 215208 4208 215260 4214
rect 215208 4150 215260 4156
rect 213932 3454 214144 3482
rect 214116 480 214144 3454
rect 215220 480 215248 4150
rect 216324 480 216352 16546
rect 217428 480 217456 16546
rect 218532 480 218560 16546
rect 219452 3194 219480 93366
rect 219532 90568 219584 90574
rect 219532 90510 219584 90516
rect 219544 16574 219572 90510
rect 223580 87848 223632 87854
rect 223580 87790 223632 87796
rect 222200 82340 222252 82346
rect 222200 82282 222252 82288
rect 220820 80912 220872 80918
rect 220820 80854 220872 80860
rect 220832 16574 220860 80854
rect 222212 16574 222240 82282
rect 223592 16574 223620 87790
rect 219544 16546 219664 16574
rect 220832 16546 221872 16574
rect 222212 16546 222976 16574
rect 223592 16546 224080 16574
rect 219440 3188 219492 3194
rect 219440 3130 219492 3136
rect 219636 480 219664 16546
rect 220728 3188 220780 3194
rect 220728 3130 220780 3136
rect 220740 480 220768 3130
rect 221844 480 221872 16546
rect 222948 480 222976 16546
rect 224052 480 224080 16546
rect 224972 3194 225000 96222
rect 226340 76764 226392 76770
rect 226340 76706 226392 76712
rect 225052 73976 225104 73982
rect 225052 73918 225104 73924
rect 225064 16574 225092 73918
rect 226352 16574 226380 76706
rect 227720 49088 227772 49094
rect 227720 49030 227772 49036
rect 227732 16574 227760 49030
rect 225064 16546 225184 16574
rect 226352 16546 227392 16574
rect 227732 16546 228496 16574
rect 224960 3188 225012 3194
rect 224960 3130 225012 3136
rect 225156 480 225184 16546
rect 226248 3188 226300 3194
rect 226248 3130 226300 3136
rect 226260 480 226288 3130
rect 227364 480 227392 16546
rect 228468 480 228496 16546
rect 229756 9654 229784 101759
rect 229848 35902 229876 109375
rect 229940 49706 229968 113183
rect 230032 74526 230060 120799
rect 230124 88330 230152 124607
rect 230386 117056 230442 117065
rect 230386 116991 230442 117000
rect 230400 116006 230428 116991
rect 230388 116000 230440 116006
rect 230388 115942 230440 115948
rect 353956 114510 353984 130319
rect 354232 128314 354260 133855
rect 354220 128308 354272 128314
rect 354220 128250 354272 128256
rect 580172 128308 580224 128314
rect 580172 128250 580224 128256
rect 580184 127673 580212 128250
rect 580170 127664 580226 127673
rect 580170 127599 580226 127608
rect 354586 126848 354642 126857
rect 354586 126783 354642 126792
rect 354494 123312 354550 123321
rect 354494 123247 354550 123256
rect 354402 119776 354458 119785
rect 354402 119711 354458 119720
rect 354310 116240 354366 116249
rect 354310 116175 354366 116184
rect 353944 114504 353996 114510
rect 353944 114446 353996 114452
rect 354218 112704 354274 112713
rect 354218 112639 354274 112648
rect 354126 109168 354182 109177
rect 354126 109103 354182 109112
rect 230386 105632 230442 105641
rect 230386 105567 230442 105576
rect 354034 105632 354090 105641
rect 354034 105567 354090 105576
rect 230400 104922 230428 105567
rect 230388 104916 230440 104922
rect 230388 104858 230440 104864
rect 353942 102096 353998 102105
rect 353942 102031 353998 102040
rect 245672 100014 246698 100042
rect 244924 97844 244976 97850
rect 244924 97786 244976 97792
rect 235264 97776 235316 97782
rect 235264 97718 235316 97724
rect 233240 92064 233292 92070
rect 233240 92006 233292 92012
rect 231860 89276 231912 89282
rect 231860 89218 231912 89224
rect 230112 88324 230164 88330
rect 230112 88266 230164 88272
rect 230480 85128 230532 85134
rect 230480 85070 230532 85076
rect 230020 74520 230072 74526
rect 230020 74462 230072 74468
rect 229928 49700 229980 49706
rect 229928 49642 229980 49648
rect 229836 35896 229888 35902
rect 229836 35838 229888 35844
rect 229744 9648 229796 9654
rect 229744 9590 229796 9596
rect 229560 9580 229612 9586
rect 229560 9522 229612 9528
rect 229572 480 229600 9522
rect 230492 3482 230520 85070
rect 230572 38004 230624 38010
rect 230572 37946 230624 37952
rect 230584 4214 230612 37946
rect 231872 16574 231900 89218
rect 233252 16574 233280 92006
rect 234620 68536 234672 68542
rect 234620 68478 234672 68484
rect 234632 16574 234660 68478
rect 235276 32434 235304 97718
rect 243544 97708 243596 97714
rect 243544 97650 243596 97656
rect 242164 97640 242216 97646
rect 242164 97582 242216 97588
rect 239404 97572 239456 97578
rect 239404 97514 239456 97520
rect 238024 97436 238076 97442
rect 238024 97378 238076 97384
rect 237380 90636 237432 90642
rect 237380 90578 237432 90584
rect 236000 86488 236052 86494
rect 236000 86430 236052 86436
rect 235264 32428 235316 32434
rect 235264 32370 235316 32376
rect 231872 16546 232912 16574
rect 233252 16546 234016 16574
rect 234632 16546 235120 16574
rect 230572 4208 230624 4214
rect 230572 4150 230624 4156
rect 231768 4208 231820 4214
rect 231768 4150 231820 4156
rect 230492 3454 230704 3482
rect 230676 480 230704 3454
rect 231780 480 231808 4150
rect 232884 480 232912 16546
rect 233988 480 234016 16546
rect 235092 480 235120 16546
rect 236012 3482 236040 86430
rect 236092 75404 236144 75410
rect 236092 75346 236144 75352
rect 236104 4214 236132 75346
rect 237392 6914 237420 90578
rect 238036 9586 238064 97378
rect 238760 94852 238812 94858
rect 238760 94794 238812 94800
rect 238024 9580 238076 9586
rect 238024 9522 238076 9528
rect 238772 6914 238800 94794
rect 239416 10402 239444 97514
rect 241520 93492 241572 93498
rect 241520 93434 241572 93440
rect 240140 83768 240192 83774
rect 240140 83710 240192 83716
rect 240152 16574 240180 83710
rect 240152 16546 240640 16574
rect 239404 10396 239456 10402
rect 239404 10338 239456 10344
rect 237392 6886 238432 6914
rect 238772 6886 239536 6914
rect 236092 4208 236144 4214
rect 236092 4150 236144 4156
rect 237288 4208 237340 4214
rect 237288 4150 237340 4156
rect 236012 3454 236224 3482
rect 236196 480 236224 3454
rect 237300 480 237328 4150
rect 238404 480 238432 6886
rect 239508 480 239536 6886
rect 240612 480 240640 16546
rect 241532 3466 241560 93434
rect 241704 15972 241756 15978
rect 241704 15914 241756 15920
rect 241428 3460 241480 3466
rect 241428 3402 241480 3408
rect 241520 3460 241572 3466
rect 241520 3402 241572 3408
rect 241440 3194 241468 3402
rect 241428 3188 241480 3194
rect 241428 3130 241480 3136
rect 241716 480 241744 15914
rect 242176 7682 242204 97582
rect 242900 61600 242952 61606
rect 242900 61542 242952 61548
rect 242912 16574 242940 61542
rect 242912 16546 243492 16574
rect 242164 7676 242216 7682
rect 242164 7618 242216 7624
rect 243464 3482 243492 16546
rect 243556 4894 243584 97650
rect 243636 96892 243688 96898
rect 243636 96834 243688 96840
rect 243648 66910 243676 96834
rect 243636 66904 243688 66910
rect 243636 66846 243688 66852
rect 244280 17400 244332 17406
rect 244280 17342 244332 17348
rect 244292 16574 244320 17342
rect 244936 17270 244964 97786
rect 244924 17264 244976 17270
rect 244924 17206 244976 17212
rect 244292 16546 245056 16574
rect 243544 4888 243596 4894
rect 243544 4830 243596 4836
rect 242808 3460 242860 3466
rect 243464 3454 243952 3482
rect 242808 3402 242860 3408
rect 242820 480 242848 3402
rect 243924 480 243952 3454
rect 245028 480 245056 16546
rect 245672 6186 245700 100014
rect 246868 96914 246896 100028
rect 246948 97912 247000 97918
rect 246948 97854 247000 97860
rect 245764 96886 246896 96914
rect 245764 6254 245792 96886
rect 246396 96824 246448 96830
rect 246396 96766 246448 96772
rect 246304 96688 246356 96694
rect 246304 96630 246356 96636
rect 245844 87916 245896 87922
rect 245844 87858 245896 87864
rect 245856 16574 245884 87858
rect 246316 37942 246344 96630
rect 246408 75206 246436 96766
rect 246960 96694 246988 97854
rect 247052 96898 247080 100028
rect 247040 96892 247092 96898
rect 247040 96834 247092 96840
rect 246948 96688 247000 96694
rect 246948 96630 247000 96636
rect 247236 93854 247264 100028
rect 247420 96914 247448 100028
rect 247604 97306 247632 100028
rect 247684 97980 247736 97986
rect 247684 97922 247736 97928
rect 247592 97300 247644 97306
rect 247592 97242 247644 97248
rect 247420 96886 247540 96914
rect 247236 93826 247448 93854
rect 246396 75200 246448 75206
rect 246396 75142 246448 75148
rect 247420 54534 247448 93826
rect 247408 54528 247460 54534
rect 247408 54470 247460 54476
rect 246304 37936 246356 37942
rect 246304 37878 246356 37884
rect 245856 16546 246160 16574
rect 245752 6248 245804 6254
rect 245752 6190 245804 6196
rect 245660 6180 245712 6186
rect 245660 6122 245712 6128
rect 246132 480 246160 16546
rect 247408 10396 247460 10402
rect 247408 10338 247460 10344
rect 247224 9036 247276 9042
rect 247224 8978 247276 8984
rect 247236 480 247264 8978
rect 247420 3074 247448 10338
rect 247512 3641 247540 96886
rect 247696 84862 247724 97922
rect 247788 96830 247816 100028
rect 247776 96824 247828 96830
rect 247776 96766 247828 96772
rect 247684 84856 247736 84862
rect 247684 84798 247736 84804
rect 247972 84194 248000 100028
rect 248156 84194 248184 100028
rect 248340 84194 248368 100028
rect 248524 97986 248552 100028
rect 248512 97980 248564 97986
rect 248512 97922 248564 97928
rect 248708 84194 248736 100028
rect 247880 84166 248000 84194
rect 248064 84166 248184 84194
rect 248248 84166 248368 84194
rect 248616 84166 248736 84194
rect 247880 31074 247908 84166
rect 247868 31068 247920 31074
rect 247868 31010 247920 31016
rect 248064 21418 248092 84166
rect 248052 21412 248104 21418
rect 248052 21354 248104 21360
rect 247498 3632 247554 3641
rect 247498 3567 247554 3576
rect 248248 3194 248276 84166
rect 248616 46238 248644 84166
rect 248892 61402 248920 100028
rect 249076 84194 249104 100028
rect 249260 97782 249288 100028
rect 249248 97776 249300 97782
rect 249248 97718 249300 97724
rect 249444 84194 249472 100028
rect 249628 84194 249656 100028
rect 249812 93854 249840 100028
rect 249996 97918 250024 100028
rect 249984 97912 250036 97918
rect 249984 97854 250036 97860
rect 250180 94518 250208 100028
rect 250168 94512 250220 94518
rect 250168 94454 250220 94460
rect 249812 93826 250024 93854
rect 248984 84166 249104 84194
rect 249352 84166 249472 84194
rect 249536 84166 249656 84194
rect 248880 61396 248932 61402
rect 248880 61338 248932 61344
rect 248604 46232 248656 46238
rect 248604 46174 248656 46180
rect 248984 3534 249012 84166
rect 249352 76566 249380 84166
rect 249340 76560 249392 76566
rect 249340 76502 249392 76508
rect 249432 4888 249484 4894
rect 249432 4830 249484 4836
rect 248972 3528 249024 3534
rect 248972 3470 249024 3476
rect 248236 3188 248288 3194
rect 248236 3130 248288 3136
rect 247420 3046 248368 3074
rect 248340 480 248368 3046
rect 249444 480 249472 4830
rect 249536 3670 249564 84166
rect 249524 3664 249576 3670
rect 249524 3606 249576 3612
rect 249996 3602 250024 93826
rect 250364 84194 250392 100028
rect 250548 84194 250576 100028
rect 250732 84194 250760 100028
rect 250916 84194 250944 100028
rect 251100 84194 251128 100028
rect 251284 84194 251312 100028
rect 250272 84166 250392 84194
rect 250456 84166 250576 84194
rect 250640 84166 250760 84194
rect 250824 84166 250944 84194
rect 251008 84166 251128 84194
rect 251192 84166 251312 84194
rect 250272 3738 250300 84166
rect 250456 3806 250484 84166
rect 250640 82142 250668 84166
rect 250628 82136 250680 82142
rect 250628 82078 250680 82084
rect 250824 36582 250852 84166
rect 250812 36576 250864 36582
rect 250812 36518 250864 36524
rect 250536 7676 250588 7682
rect 250536 7618 250588 7624
rect 250444 3800 250496 3806
rect 250444 3742 250496 3748
rect 250260 3732 250312 3738
rect 250260 3674 250312 3680
rect 249984 3596 250036 3602
rect 249984 3538 250036 3544
rect 250548 480 250576 7618
rect 251008 3874 251036 84166
rect 251192 72486 251220 84166
rect 251180 72480 251232 72486
rect 251180 72422 251232 72428
rect 251468 33794 251496 100028
rect 251652 84194 251680 100028
rect 251836 84194 251864 100028
rect 252020 84194 252048 100028
rect 252204 84194 252232 100028
rect 252388 84194 252416 100028
rect 251560 84166 251680 84194
rect 251744 84166 251864 84194
rect 251928 84166 252048 84194
rect 252112 84166 252232 84194
rect 252296 84166 252416 84194
rect 251456 33788 251508 33794
rect 251456 33730 251508 33736
rect 251560 3942 251588 84166
rect 251744 64190 251772 84166
rect 251732 64184 251784 64190
rect 251732 64126 251784 64132
rect 251928 10334 251956 84166
rect 251916 10328 251968 10334
rect 251916 10270 251968 10276
rect 251640 7744 251692 7750
rect 251640 7686 251692 7692
rect 251548 3936 251600 3942
rect 251548 3878 251600 3884
rect 250996 3868 251048 3874
rect 250996 3810 251048 3816
rect 251652 480 251680 7686
rect 252112 4010 252140 84166
rect 252296 55894 252324 84166
rect 252572 83502 252600 100028
rect 252756 84194 252784 100028
rect 252940 96830 252968 100028
rect 253124 96914 253152 100028
rect 253032 96886 253152 96914
rect 252928 96824 252980 96830
rect 252928 96766 252980 96772
rect 252664 84166 252784 84194
rect 252560 83496 252612 83502
rect 252560 83438 252612 83444
rect 252284 55888 252336 55894
rect 252284 55830 252336 55836
rect 252664 4078 252692 84166
rect 253032 68338 253060 96886
rect 253112 96824 253164 96830
rect 253112 96766 253164 96772
rect 253124 93158 253152 96766
rect 253112 93152 253164 93158
rect 253112 93094 253164 93100
rect 253308 84194 253336 100028
rect 253492 84194 253520 100028
rect 253676 84194 253704 100028
rect 253860 84194 253888 100028
rect 254044 93226 254072 100028
rect 254032 93220 254084 93226
rect 254032 93162 254084 93168
rect 254228 84194 254256 100028
rect 253216 84166 253336 84194
rect 253400 84166 253520 84194
rect 253584 84166 253704 84194
rect 253768 84166 253888 84194
rect 254136 84166 254256 84194
rect 253020 68332 253072 68338
rect 253020 68274 253072 68280
rect 252744 6180 252796 6186
rect 252744 6122 252796 6128
rect 252652 4072 252704 4078
rect 252652 4014 252704 4020
rect 252100 4004 252152 4010
rect 252100 3946 252152 3952
rect 252756 480 252784 6122
rect 253216 4146 253244 84166
rect 253400 65550 253428 84166
rect 253388 65544 253440 65550
rect 253388 65486 253440 65492
rect 253584 22778 253612 84166
rect 253572 22772 253624 22778
rect 253572 22714 253624 22720
rect 253204 4140 253256 4146
rect 253204 4082 253256 4088
rect 253768 3398 253796 84166
rect 254136 29646 254164 84166
rect 254124 29640 254176 29646
rect 254124 29582 254176 29588
rect 254412 7614 254440 100028
rect 254596 94586 254624 100028
rect 254584 94580 254636 94586
rect 254584 94522 254636 94528
rect 254780 84194 254808 100028
rect 254964 84194 254992 100028
rect 255148 84194 255176 100028
rect 255332 94450 255360 100028
rect 255516 96914 255544 100028
rect 255700 97850 255728 100028
rect 255688 97844 255740 97850
rect 255688 97786 255740 97792
rect 255424 96886 255544 96914
rect 255320 94444 255372 94450
rect 255320 94386 255372 94392
rect 254688 84166 254808 84194
rect 254872 84166 254992 84194
rect 255056 84166 255176 84194
rect 254688 51746 254716 84166
rect 254676 51740 254728 51746
rect 254676 51682 254728 51688
rect 254872 11762 254900 84166
rect 255056 83570 255084 84166
rect 255044 83564 255096 83570
rect 255044 83506 255096 83512
rect 255424 19990 255452 96886
rect 255504 94444 255556 94450
rect 255504 94386 255556 94392
rect 255516 53106 255544 94386
rect 255504 53100 255556 53106
rect 255504 53042 255556 53048
rect 255884 50386 255912 100028
rect 255964 97164 256016 97170
rect 255964 97106 256016 97112
rect 255976 86290 256004 97106
rect 255964 86284 256016 86290
rect 255964 86226 256016 86232
rect 255872 50380 255924 50386
rect 255872 50322 255924 50328
rect 255412 19984 255464 19990
rect 255412 19926 255464 19932
rect 256068 18630 256096 100028
rect 256252 95946 256280 100028
rect 256240 95940 256292 95946
rect 256240 95882 256292 95888
rect 256436 84194 256464 100028
rect 256620 84194 256648 100028
rect 256804 89010 256832 100028
rect 256988 93854 257016 100028
rect 257172 96014 257200 100028
rect 257356 96914 257384 100028
rect 257436 97028 257488 97034
rect 257436 96970 257488 96976
rect 257264 96886 257384 96914
rect 257160 96008 257212 96014
rect 257160 95950 257212 95956
rect 256988 93826 257200 93854
rect 256792 89004 256844 89010
rect 256792 88946 256844 88952
rect 256344 84166 256464 84194
rect 256528 84166 256648 84194
rect 256344 28286 256372 84166
rect 256528 77994 256556 84166
rect 256516 77988 256568 77994
rect 256516 77930 256568 77936
rect 256332 28280 256384 28286
rect 256332 28222 256384 28228
rect 257172 26926 257200 93826
rect 257264 76634 257292 96886
rect 257344 96688 257396 96694
rect 257344 96630 257396 96636
rect 257252 76628 257304 76634
rect 257252 76570 257304 76576
rect 257160 26920 257212 26926
rect 257160 26862 257212 26868
rect 257356 24138 257384 96630
rect 257448 90370 257476 96970
rect 257436 90364 257488 90370
rect 257436 90306 257488 90312
rect 257540 39370 257568 100028
rect 257724 84194 257752 100028
rect 257908 84194 257936 100028
rect 258092 96694 258120 100028
rect 258080 96688 258132 96694
rect 258080 96630 258132 96636
rect 258276 84930 258304 100028
rect 258460 97170 258488 100028
rect 258448 97164 258500 97170
rect 258448 97106 258500 97112
rect 258264 84924 258316 84930
rect 258264 84866 258316 84872
rect 257632 84166 257752 84194
rect 257816 84166 257936 84194
rect 257528 39364 257580 39370
rect 257528 39306 257580 39312
rect 257344 24132 257396 24138
rect 257344 24074 257396 24080
rect 256056 18624 256108 18630
rect 256056 18566 256108 18572
rect 254860 11756 254912 11762
rect 254860 11698 254912 11704
rect 257160 10328 257212 10334
rect 257160 10270 257212 10276
rect 254400 7608 254452 7614
rect 254400 7550 254452 7556
rect 253848 6384 253900 6390
rect 253848 6326 253900 6332
rect 253756 3392 253808 3398
rect 253756 3334 253808 3340
rect 253860 480 253888 6326
rect 256056 5024 256108 5030
rect 256056 4966 256108 4972
rect 254952 4956 255004 4962
rect 254952 4898 255004 4904
rect 254964 480 254992 4898
rect 256068 480 256096 4966
rect 257172 480 257200 10270
rect 257632 4826 257660 84166
rect 257816 68406 257844 84166
rect 258644 73846 258672 100028
rect 258828 84194 258856 100028
rect 259012 97034 259040 100028
rect 259000 97028 259052 97034
rect 259000 96970 259052 96976
rect 259196 84194 259224 100028
rect 259380 84194 259408 100028
rect 259564 96914 259592 100028
rect 258736 84166 258856 84194
rect 259104 84166 259224 84194
rect 259288 84166 259408 84194
rect 259472 96886 259592 96914
rect 258632 73840 258684 73846
rect 258632 73782 258684 73788
rect 257804 68400 257856 68406
rect 257804 68342 257856 68348
rect 258736 32502 258764 84166
rect 259104 47598 259132 84166
rect 259092 47592 259144 47598
rect 259092 47534 259144 47540
rect 258724 32496 258776 32502
rect 258724 32438 258776 32444
rect 259288 31142 259316 84166
rect 259472 79354 259500 96886
rect 259748 84194 259776 100028
rect 259932 89078 259960 100028
rect 260116 96914 260144 100028
rect 260024 96886 260144 96914
rect 259920 89072 259972 89078
rect 259920 89014 259972 89020
rect 259564 84166 259776 84194
rect 259460 79348 259512 79354
rect 259460 79290 259512 79296
rect 259276 31136 259328 31142
rect 259276 31078 259328 31084
rect 259564 25566 259592 84166
rect 260024 78062 260052 96886
rect 260104 96756 260156 96762
rect 260104 96698 260156 96704
rect 260012 78056 260064 78062
rect 260012 77998 260064 78004
rect 260116 69698 260144 96698
rect 260300 84194 260328 100028
rect 260484 84194 260512 100028
rect 260668 84194 260696 100028
rect 260852 96914 260880 100028
rect 261036 97034 261064 100028
rect 261024 97028 261076 97034
rect 261024 96970 261076 96976
rect 260852 96886 261064 96914
rect 260932 96824 260984 96830
rect 260932 96766 260984 96772
rect 260208 84166 260328 84194
rect 260392 84166 260512 84194
rect 260576 84166 260696 84194
rect 260104 69692 260156 69698
rect 260104 69634 260156 69640
rect 259552 25560 259604 25566
rect 259552 25502 259604 25508
rect 260208 15910 260236 84166
rect 260392 29714 260420 84166
rect 260576 62830 260604 84166
rect 260564 62824 260616 62830
rect 260564 62766 260616 62772
rect 260944 44878 260972 96766
rect 261036 75274 261064 96886
rect 261220 91798 261248 100028
rect 261404 96830 261432 100028
rect 261484 97028 261536 97034
rect 261484 96970 261536 96976
rect 261392 96824 261444 96830
rect 261392 96766 261444 96772
rect 261208 91792 261260 91798
rect 261208 91734 261260 91740
rect 261024 75268 261076 75274
rect 261024 75210 261076 75216
rect 260932 44872 260984 44878
rect 260932 44814 260984 44820
rect 260380 29708 260432 29714
rect 260380 29650 260432 29656
rect 260196 15904 260248 15910
rect 260196 15846 260248 15852
rect 261496 9178 261524 96970
rect 261588 17338 261616 100028
rect 261772 84194 261800 100028
rect 261956 84194 261984 100028
rect 262140 84194 262168 100028
rect 262324 96762 262352 100028
rect 262312 96756 262364 96762
rect 262312 96698 262364 96704
rect 261680 84166 261800 84194
rect 261864 84166 261984 84194
rect 262048 84166 262168 84194
rect 261680 71058 261708 84166
rect 261668 71052 261720 71058
rect 261668 70994 261720 71000
rect 261864 40730 261892 84166
rect 261852 40724 261904 40730
rect 261852 40666 261904 40672
rect 262048 28354 262076 84166
rect 262508 66978 262536 100028
rect 262496 66972 262548 66978
rect 262496 66914 262548 66920
rect 262036 28348 262088 28354
rect 262036 28290 262088 28296
rect 262692 26994 262720 100028
rect 262876 87650 262904 100028
rect 262864 87644 262916 87650
rect 262864 87586 262916 87592
rect 263060 84194 263088 100028
rect 263244 84194 263272 100028
rect 263428 84194 263456 100028
rect 263612 96914 263640 100028
rect 263796 97374 263824 100028
rect 263784 97368 263836 97374
rect 263784 97310 263836 97316
rect 263612 96886 263824 96914
rect 263692 96824 263744 96830
rect 263692 96766 263744 96772
rect 262968 84166 263088 84194
rect 263152 84166 263272 84194
rect 263336 84166 263456 84194
rect 262968 42090 262996 84166
rect 262956 42084 263008 42090
rect 262956 42026 263008 42032
rect 262680 26988 262732 26994
rect 262680 26930 262732 26936
rect 263152 24206 263180 84166
rect 263336 80714 263364 84166
rect 263324 80708 263376 80714
rect 263324 80650 263376 80656
rect 263140 24200 263192 24206
rect 263140 24142 263192 24148
rect 261576 17332 261628 17338
rect 261576 17274 261628 17280
rect 263704 14482 263732 96766
rect 263796 43450 263824 96886
rect 263980 84194 264008 100028
rect 264164 96830 264192 100028
rect 264244 96892 264296 96898
rect 264244 96834 264296 96840
rect 264152 96824 264204 96830
rect 264152 96766 264204 96772
rect 264256 86358 264284 96834
rect 264244 86352 264296 86358
rect 264244 86294 264296 86300
rect 263888 84166 264008 84194
rect 263888 61470 263916 84166
rect 263876 61464 263928 61470
rect 263876 61406 263928 61412
rect 263784 43444 263836 43450
rect 263784 43386 263836 43392
rect 264348 25634 264376 100028
rect 264532 84194 264560 100028
rect 264716 84194 264744 100028
rect 264900 97510 264928 100028
rect 264888 97504 264940 97510
rect 264888 97446 264940 97452
rect 264980 97232 265032 97238
rect 264980 97174 265032 97180
rect 264992 94654 265020 97174
rect 264980 94648 265032 94654
rect 264980 94590 265032 94596
rect 264440 84166 264560 84194
rect 264624 84166 264744 84194
rect 264440 60042 264468 84166
rect 264428 60036 264480 60042
rect 264428 59978 264480 59984
rect 264336 25628 264388 25634
rect 264336 25570 264388 25576
rect 263692 14476 263744 14482
rect 263692 14418 263744 14424
rect 264624 13122 264652 84166
rect 265084 58682 265112 100028
rect 265164 96960 265216 96966
rect 265164 96902 265216 96908
rect 265072 58676 265124 58682
rect 265072 58618 265124 58624
rect 265176 57254 265204 96902
rect 265164 57248 265216 57254
rect 265164 57190 265216 57196
rect 265268 49026 265296 100028
rect 265452 93854 265480 100028
rect 265636 96966 265664 100028
rect 265624 96960 265676 96966
rect 265624 96902 265676 96908
rect 265624 96756 265676 96762
rect 265624 96698 265676 96704
rect 265452 93826 265572 93854
rect 265256 49020 265308 49026
rect 265256 48962 265308 48968
rect 264612 13116 264664 13122
rect 264612 13058 264664 13064
rect 263784 11756 263836 11762
rect 263784 11698 263836 11704
rect 261484 9172 261536 9178
rect 261484 9114 261536 9120
rect 260472 9104 260524 9110
rect 260472 9046 260524 9052
rect 258264 6248 258316 6254
rect 258264 6190 258316 6196
rect 257620 4820 257672 4826
rect 257620 4762 257672 4768
rect 258276 480 258304 6190
rect 259368 4820 259420 4826
rect 259368 4762 259420 4768
rect 259380 480 259408 4762
rect 260484 480 260512 9046
rect 261576 8968 261628 8974
rect 261576 8910 261628 8916
rect 261588 480 261616 8910
rect 262680 6316 262732 6322
rect 262680 6258 262732 6264
rect 262692 480 262720 6258
rect 263796 480 263824 11698
rect 264888 3460 264940 3466
rect 264888 3402 264940 3408
rect 264900 480 264928 3402
rect 265544 3330 265572 93826
rect 265636 80782 265664 96698
rect 265624 80776 265676 80782
rect 265624 80718 265676 80724
rect 265820 35222 265848 100028
rect 266004 84194 266032 100028
rect 266188 97714 266216 100028
rect 266176 97708 266228 97714
rect 266176 97650 266228 97656
rect 266372 89146 266400 100028
rect 266360 89140 266412 89146
rect 266360 89082 266412 89088
rect 266556 84194 266584 100028
rect 266740 96898 266768 100028
rect 266728 96892 266780 96898
rect 266728 96834 266780 96840
rect 266924 84194 266952 100028
rect 267108 84194 267136 100028
rect 267292 96762 267320 100028
rect 267280 96756 267332 96762
rect 267280 96698 267332 96704
rect 267476 84194 267504 100028
rect 267660 84194 267688 100028
rect 267844 84194 267872 100028
rect 265912 84166 266032 84194
rect 266464 84166 266584 84194
rect 266832 84166 266952 84194
rect 267016 84166 267136 84194
rect 267384 84166 267504 84194
rect 267568 84166 267688 84194
rect 267752 84166 267872 84194
rect 265808 35216 265860 35222
rect 265808 35158 265860 35164
rect 265532 3324 265584 3330
rect 265532 3266 265584 3272
rect 265912 3262 265940 84166
rect 266464 82210 266492 84166
rect 266452 82204 266504 82210
rect 266452 82146 266504 82152
rect 266832 65618 266860 84166
rect 266820 65612 266872 65618
rect 266820 65554 266872 65560
rect 266452 63028 266504 63034
rect 266452 62970 266504 62976
rect 266464 16574 266492 62970
rect 267016 43518 267044 84166
rect 267384 62898 267412 84166
rect 267372 62892 267424 62898
rect 267372 62834 267424 62840
rect 267004 43512 267056 43518
rect 267004 43454 267056 43460
rect 267568 36650 267596 84166
rect 267752 79422 267780 84166
rect 267740 79416 267792 79422
rect 267740 79358 267792 79364
rect 268028 60110 268056 100028
rect 268212 93854 268240 100028
rect 268212 93826 268332 93854
rect 268016 60104 268068 60110
rect 268016 60046 268068 60052
rect 267556 36644 267608 36650
rect 267556 36586 267608 36592
rect 268304 18698 268332 93826
rect 268396 84998 268424 100028
rect 268384 84992 268436 84998
rect 268384 84934 268436 84940
rect 268580 84194 268608 100028
rect 268764 84194 268792 100028
rect 268948 84194 268976 100028
rect 269132 95266 269160 100028
rect 269316 96914 269344 100028
rect 269224 96886 269344 96914
rect 269120 95260 269172 95266
rect 269120 95202 269172 95208
rect 268488 84166 268608 84194
rect 268672 84166 268792 84194
rect 268856 84166 268976 84194
rect 268488 58750 268516 84166
rect 268476 58744 268528 58750
rect 268476 58686 268528 58692
rect 268672 33862 268700 84166
rect 268856 78130 268884 84166
rect 268844 78124 268896 78130
rect 268844 78066 268896 78072
rect 268660 33856 268712 33862
rect 268660 33798 268712 33804
rect 269224 20058 269252 96886
rect 269396 96620 269448 96626
rect 269396 96562 269448 96568
rect 269408 96150 269436 96562
rect 269500 96150 269528 100028
rect 269684 96914 269712 100028
rect 269592 96886 269712 96914
rect 269396 96144 269448 96150
rect 269396 96086 269448 96092
rect 269488 96144 269540 96150
rect 269488 96086 269540 96092
rect 269304 95260 269356 95266
rect 269304 95202 269356 95208
rect 269316 72554 269344 95202
rect 269304 72548 269356 72554
rect 269304 72490 269356 72496
rect 269592 57322 269620 96886
rect 269672 96144 269724 96150
rect 269672 96086 269724 96092
rect 269684 91866 269712 96086
rect 269672 91860 269724 91866
rect 269672 91802 269724 91808
rect 269868 84194 269896 100028
rect 270052 84194 270080 100028
rect 270236 84194 270264 100028
rect 270420 84194 270448 100028
rect 270604 84194 270632 100028
rect 269776 84166 269896 84194
rect 269960 84166 270080 84194
rect 270144 84166 270264 84194
rect 270328 84166 270448 84194
rect 270512 84166 270632 84194
rect 269580 57316 269632 57322
rect 269580 57258 269632 57264
rect 269212 20052 269264 20058
rect 269212 19994 269264 20000
rect 268292 18692 268344 18698
rect 268292 18634 268344 18640
rect 266464 16546 267136 16574
rect 265992 7608 266044 7614
rect 265992 7550 266044 7556
rect 265900 3256 265952 3262
rect 265900 3198 265952 3204
rect 266004 480 266032 7550
rect 267108 480 267136 16546
rect 269776 11830 269804 84166
rect 269960 83638 269988 84166
rect 269948 83632 270000 83638
rect 269948 83574 270000 83580
rect 270144 55962 270172 84166
rect 270328 64258 270356 84166
rect 270512 76702 270540 84166
rect 270500 76696 270552 76702
rect 270500 76638 270552 76644
rect 270316 64252 270368 64258
rect 270316 64194 270368 64200
rect 270132 55956 270184 55962
rect 270132 55898 270184 55904
rect 270788 54602 270816 100028
rect 270776 54596 270828 54602
rect 270776 54538 270828 54544
rect 270972 21486 271000 100028
rect 271156 96914 271184 100028
rect 271064 96886 271184 96914
rect 271064 82278 271092 96886
rect 271144 96824 271196 96830
rect 271144 96766 271196 96772
rect 271052 82272 271104 82278
rect 271052 82214 271104 82220
rect 271156 75342 271184 96766
rect 271340 84194 271368 100028
rect 271524 84194 271552 100028
rect 271708 96082 271736 100028
rect 271892 96830 271920 100028
rect 271880 96824 271932 96830
rect 271880 96766 271932 96772
rect 271696 96076 271748 96082
rect 271696 96018 271748 96024
rect 271248 84166 271368 84194
rect 271432 84166 271552 84194
rect 271144 75336 271196 75342
rect 271144 75278 271196 75284
rect 271248 53174 271276 84166
rect 271236 53168 271288 53174
rect 271236 53110 271288 53116
rect 271432 22846 271460 84166
rect 272076 61538 272104 100028
rect 272260 97646 272288 100028
rect 272248 97640 272300 97646
rect 272248 97582 272300 97588
rect 272444 90438 272472 100028
rect 272524 96892 272576 96898
rect 272524 96834 272576 96840
rect 272432 90432 272484 90438
rect 272432 90374 272484 90380
rect 272536 87718 272564 96834
rect 272524 87712 272576 87718
rect 272524 87654 272576 87660
rect 272064 61532 272116 61538
rect 272064 61474 272116 61480
rect 272628 51814 272656 100028
rect 272812 97238 272840 100028
rect 272800 97232 272852 97238
rect 272800 97174 272852 97180
rect 272996 84194 273024 100028
rect 273180 84194 273208 100028
rect 273364 93294 273392 100028
rect 273352 93288 273404 93294
rect 273352 93230 273404 93236
rect 272904 84166 273024 84194
rect 273088 84166 273208 84194
rect 272904 72622 272932 84166
rect 272892 72616 272944 72622
rect 272892 72558 272944 72564
rect 272616 51808 272668 51814
rect 272616 51750 272668 51756
rect 273088 50454 273116 84166
rect 273548 71126 273576 100028
rect 273628 96960 273680 96966
rect 273628 96902 273680 96908
rect 273536 71120 273588 71126
rect 273536 71062 273588 71068
rect 273260 71052 273312 71058
rect 273260 70994 273312 71000
rect 273076 50448 273128 50454
rect 273076 50390 273128 50396
rect 271420 22840 271472 22846
rect 271420 22782 271472 22788
rect 270960 21480 271012 21486
rect 270960 21422 271012 21428
rect 273272 16574 273300 70994
rect 273640 69766 273668 96902
rect 273628 69760 273680 69766
rect 273628 69702 273680 69708
rect 273732 47666 273760 100028
rect 273916 96914 273944 100028
rect 273996 97300 274048 97306
rect 273996 97242 274048 97248
rect 273824 96886 273944 96914
rect 273824 91934 273852 96886
rect 274008 95554 274036 97242
rect 274100 96966 274128 100028
rect 274180 97028 274232 97034
rect 274180 96970 274232 96976
rect 274088 96960 274140 96966
rect 274088 96902 274140 96908
rect 274088 96756 274140 96762
rect 274088 96698 274140 96704
rect 273916 95526 274036 95554
rect 273812 91928 273864 91934
rect 273812 91870 273864 91876
rect 273720 47660 273772 47666
rect 273720 47602 273772 47608
rect 273272 16546 273760 16574
rect 269764 11824 269816 11830
rect 269764 11766 269816 11772
rect 270408 6452 270460 6458
rect 270408 6394 270460 6400
rect 269304 5092 269356 5098
rect 269304 5034 269356 5040
rect 268200 3528 268252 3534
rect 268200 3470 268252 3476
rect 268212 480 268240 3470
rect 269316 480 269344 5034
rect 270420 480 270448 6394
rect 272616 5160 272668 5166
rect 272616 5102 272668 5108
rect 271512 3596 271564 3602
rect 271512 3538 271564 3544
rect 271524 480 271552 3538
rect 272628 480 272656 5102
rect 273732 480 273760 16546
rect 273916 5030 273944 95526
rect 273996 95464 274048 95470
rect 273996 95406 274048 95412
rect 274008 85066 274036 95406
rect 274100 90506 274128 96698
rect 274192 95470 274220 96970
rect 274180 95464 274232 95470
rect 274180 95406 274232 95412
rect 274088 90500 274140 90506
rect 274088 90442 274140 90448
rect 273996 85060 274048 85066
rect 273996 85002 274048 85008
rect 274284 84194 274312 100028
rect 274468 97578 274496 100028
rect 274456 97572 274508 97578
rect 274456 97514 274508 97520
rect 274652 93854 274680 100028
rect 274836 96898 274864 100028
rect 274824 96892 274876 96898
rect 274824 96834 274876 96840
rect 275020 96762 275048 100028
rect 275100 96960 275152 96966
rect 275100 96902 275152 96908
rect 275008 96756 275060 96762
rect 275008 96698 275060 96704
rect 274652 93826 274956 93854
rect 274192 84166 274312 84194
rect 274192 46306 274220 84166
rect 274928 68474 274956 93826
rect 274916 68468 274968 68474
rect 274916 68410 274968 68416
rect 274180 46300 274232 46306
rect 274180 46242 274232 46248
rect 275112 44946 275140 96902
rect 275204 80850 275232 100028
rect 275284 97504 275336 97510
rect 275284 97446 275336 97452
rect 275192 80844 275244 80850
rect 275192 80786 275244 80792
rect 275100 44940 275152 44946
rect 275100 44882 275152 44888
rect 275296 6390 275324 97446
rect 275388 96966 275416 100028
rect 275376 96960 275428 96966
rect 275376 96902 275428 96908
rect 275572 89214 275600 100028
rect 275560 89208 275612 89214
rect 275560 89150 275612 89156
rect 275756 84194 275784 100028
rect 275940 84194 275968 100028
rect 276124 96694 276152 100028
rect 276112 96688 276164 96694
rect 276112 96630 276164 96636
rect 276308 86426 276336 100028
rect 276296 86420 276348 86426
rect 276296 86362 276348 86368
rect 276492 84194 276520 100028
rect 276676 97322 276704 100028
rect 276756 97912 276808 97918
rect 276756 97854 276808 97860
rect 276584 97294 276704 97322
rect 276584 94722 276612 97294
rect 276664 96756 276716 96762
rect 276664 96698 276716 96704
rect 276572 94716 276624 94722
rect 276572 94658 276624 94664
rect 275664 84166 275784 84194
rect 275848 84166 275968 84194
rect 276400 84166 276520 84194
rect 275664 67046 275692 84166
rect 275652 67040 275704 67046
rect 275652 66982 275704 66988
rect 275848 13190 275876 84166
rect 276020 73840 276072 73846
rect 276020 73782 276072 73788
rect 276032 16574 276060 73782
rect 276400 71194 276428 84166
rect 276388 71188 276440 71194
rect 276388 71130 276440 71136
rect 276676 42158 276704 96698
rect 276768 93362 276796 97854
rect 276756 93356 276808 93362
rect 276756 93298 276808 93304
rect 276860 73914 276888 100028
rect 277044 84194 277072 100028
rect 277228 97034 277256 100028
rect 277216 97028 277268 97034
rect 277216 96970 277268 96976
rect 277412 93854 277440 100028
rect 277596 96762 277624 100028
rect 277780 97918 277808 100028
rect 277768 97912 277820 97918
rect 277768 97854 277820 97860
rect 277584 96756 277636 96762
rect 277584 96698 277636 96704
rect 277860 95736 277912 95742
rect 277860 95678 277912 95684
rect 277412 93826 277716 93854
rect 276952 84166 277072 84194
rect 276848 73908 276900 73914
rect 276848 73850 276900 73856
rect 276952 69834 276980 84166
rect 277688 79490 277716 93826
rect 277676 79484 277728 79490
rect 277676 79426 277728 79432
rect 276940 69828 276992 69834
rect 276940 69770 276992 69776
rect 276664 42152 276716 42158
rect 276664 42094 276716 42100
rect 276032 16546 277072 16574
rect 275836 13184 275888 13190
rect 275836 13126 275888 13132
rect 275928 6928 275980 6934
rect 275928 6870 275980 6876
rect 275284 6384 275336 6390
rect 275284 6326 275336 6332
rect 273904 5024 273956 5030
rect 273904 4966 273956 4972
rect 274824 3664 274876 3670
rect 274824 3606 274876 3612
rect 274836 480 274864 3606
rect 275940 480 275968 6870
rect 277044 480 277072 16546
rect 277872 14550 277900 95678
rect 277964 78198 277992 100028
rect 278044 97368 278096 97374
rect 278044 97310 278096 97316
rect 277952 78192 278004 78198
rect 277952 78134 278004 78140
rect 277860 14544 277912 14550
rect 277860 14486 277912 14492
rect 278056 6458 278084 97310
rect 278148 95742 278176 100028
rect 278228 97300 278280 97306
rect 278228 97242 278280 97248
rect 278136 95736 278188 95742
rect 278136 95678 278188 95684
rect 278240 94790 278268 97242
rect 278228 94784 278280 94790
rect 278228 94726 278280 94732
rect 278332 87786 278360 100028
rect 278412 97640 278464 97646
rect 278412 97582 278464 97588
rect 278424 96286 278452 97582
rect 278412 96280 278464 96286
rect 278412 96222 278464 96228
rect 278320 87780 278372 87786
rect 278320 87722 278372 87728
rect 278516 84194 278544 100028
rect 278700 84194 278728 100028
rect 278884 92002 278912 100028
rect 279068 97306 279096 100028
rect 279056 97300 279108 97306
rect 279056 97242 279108 97248
rect 278872 91996 278924 92002
rect 278872 91938 278924 91944
rect 279252 84194 279280 100028
rect 279436 96948 279464 100028
rect 279620 98138 279648 100028
rect 278424 84166 278544 84194
rect 278608 84166 278728 84194
rect 279160 84166 279280 84194
rect 279344 96920 279464 96948
rect 279528 98110 279648 98138
rect 278424 64326 278452 84166
rect 278412 64320 278464 64326
rect 278412 64262 278464 64268
rect 278608 40798 278636 84166
rect 279160 65686 279188 84166
rect 279344 83706 279372 96920
rect 279424 96688 279476 96694
rect 279424 96630 279476 96636
rect 279436 95690 279464 96630
rect 279528 96218 279556 98110
rect 279608 96960 279660 96966
rect 279608 96902 279660 96908
rect 279516 96212 279568 96218
rect 279516 96154 279568 96160
rect 279436 95662 279556 95690
rect 279424 95600 279476 95606
rect 279424 95542 279476 95548
rect 279332 83700 279384 83706
rect 279332 83642 279384 83648
rect 279148 65680 279200 65686
rect 279148 65622 279200 65628
rect 278596 40792 278648 40798
rect 278596 40734 278648 40740
rect 279240 9172 279292 9178
rect 279240 9114 279292 9120
rect 278044 6452 278096 6458
rect 278044 6394 278096 6400
rect 278136 3732 278188 3738
rect 278136 3674 278188 3680
rect 278148 480 278176 3674
rect 279252 480 279280 9114
rect 279436 4826 279464 95542
rect 279528 6934 279556 95662
rect 279620 82346 279648 96902
rect 279700 96892 279752 96898
rect 279700 96834 279752 96840
rect 279712 95606 279740 96834
rect 279700 95600 279752 95606
rect 279700 95542 279752 95548
rect 279804 84194 279832 100028
rect 279884 97572 279936 97578
rect 279884 97514 279936 97520
rect 279896 96694 279924 97514
rect 279884 96688 279936 96694
rect 279884 96630 279936 96636
rect 279988 90574 280016 100028
rect 280172 93430 280200 100028
rect 280160 93424 280212 93430
rect 280160 93366 280212 93372
rect 279976 90568 280028 90574
rect 279976 90510 280028 90516
rect 279712 84166 279832 84194
rect 279608 82340 279660 82346
rect 279608 82282 279660 82288
rect 279712 39438 279740 84166
rect 280356 80918 280384 100028
rect 280540 96966 280568 100028
rect 280528 96960 280580 96966
rect 280528 96902 280580 96908
rect 280724 87854 280752 100028
rect 280712 87848 280764 87854
rect 280712 87790 280764 87796
rect 280908 84194 280936 100028
rect 281092 97646 281120 100028
rect 281080 97640 281132 97646
rect 281080 97582 281132 97588
rect 281276 84194 281304 100028
rect 281460 84194 281488 100028
rect 281644 97442 281672 100028
rect 281632 97436 281684 97442
rect 281632 97378 281684 97384
rect 281540 97232 281592 97238
rect 281540 97174 281592 97180
rect 281552 94858 281580 97174
rect 281632 95192 281684 95198
rect 281632 95134 281684 95140
rect 281540 94852 281592 94858
rect 281540 94794 281592 94800
rect 281644 92070 281672 95134
rect 281632 92064 281684 92070
rect 281632 92006 281684 92012
rect 281828 85134 281856 100028
rect 281816 85128 281868 85134
rect 281816 85070 281868 85076
rect 282012 84194 282040 100028
rect 282196 96948 282224 100028
rect 282276 97844 282328 97850
rect 282276 97786 282328 97792
rect 282104 96920 282224 96948
rect 282104 89282 282132 96920
rect 282184 96824 282236 96830
rect 282184 96766 282236 96772
rect 282092 89276 282144 89282
rect 282092 89218 282144 89224
rect 280816 84166 280936 84194
rect 281184 84166 281304 84194
rect 281368 84166 281488 84194
rect 281920 84166 282040 84194
rect 280344 80912 280396 80918
rect 280344 80854 280396 80860
rect 280816 73982 280844 84166
rect 281184 76770 281212 84166
rect 281172 76764 281224 76770
rect 281172 76706 281224 76712
rect 280804 73976 280856 73982
rect 280804 73918 280856 73924
rect 281368 49094 281396 84166
rect 281356 49088 281408 49094
rect 281356 49030 281408 49036
rect 279700 39432 279752 39438
rect 279700 39374 279752 39380
rect 281920 38010 281948 84166
rect 281908 38004 281960 38010
rect 281908 37946 281960 37952
rect 279516 6928 279568 6934
rect 279516 6870 279568 6876
rect 280344 5568 280396 5574
rect 280344 5510 280396 5516
rect 279424 4820 279476 4826
rect 279424 4762 279476 4768
rect 280356 480 280384 5510
rect 282196 4894 282224 96766
rect 282288 5166 282316 97786
rect 282380 95198 282408 100028
rect 282368 95192 282420 95198
rect 282368 95134 282420 95140
rect 282564 84194 282592 100028
rect 282748 86494 282776 100028
rect 282932 93854 282960 100028
rect 283116 96694 283144 100028
rect 283300 97238 283328 100028
rect 283288 97232 283340 97238
rect 283288 97174 283340 97180
rect 283484 96948 283512 100028
rect 283208 96920 283512 96948
rect 283104 96688 283156 96694
rect 283104 96630 283156 96636
rect 282932 93826 283052 93854
rect 282736 86488 282788 86494
rect 282736 86430 282788 86436
rect 282472 84166 282592 84194
rect 282472 68542 282500 84166
rect 283024 75410 283052 93826
rect 283208 83774 283236 96920
rect 283668 96778 283696 100028
rect 283392 96750 283696 96778
rect 283196 83768 283248 83774
rect 283196 83710 283248 83716
rect 283012 75404 283064 75410
rect 283012 75346 283064 75352
rect 282460 68536 282512 68542
rect 282460 68478 282512 68484
rect 283392 15978 283420 96750
rect 283472 96688 283524 96694
rect 283472 96630 283524 96636
rect 283564 96688 283616 96694
rect 283564 96630 283616 96636
rect 283656 96688 283708 96694
rect 283656 96630 283708 96636
rect 283484 90642 283512 96630
rect 283472 90636 283524 90642
rect 283472 90578 283524 90584
rect 283380 15972 283432 15978
rect 283380 15914 283432 15920
rect 282276 5160 282328 5166
rect 282276 5102 282328 5108
rect 283576 4962 283604 96630
rect 283668 9042 283696 96630
rect 283852 93498 283880 100028
rect 283840 93492 283892 93498
rect 283840 93434 283892 93440
rect 284036 84194 284064 100028
rect 284220 84194 284248 100028
rect 284404 87922 284432 100028
rect 284588 96694 284616 100028
rect 284576 96688 284628 96694
rect 284576 96630 284628 96636
rect 284392 87916 284444 87922
rect 284392 87858 284444 87864
rect 284772 84194 284800 100028
rect 284956 98002 284984 100028
rect 284864 97974 284984 98002
rect 284864 96830 284892 97974
rect 284944 97912 284996 97918
rect 284944 97854 284996 97860
rect 284852 96824 284904 96830
rect 284852 96766 284904 96772
rect 283944 84166 284064 84194
rect 284128 84166 284248 84194
rect 284680 84166 284800 84194
rect 283944 61606 283972 84166
rect 283932 61600 283984 61606
rect 283932 61542 283984 61548
rect 284128 17406 284156 84166
rect 284116 17400 284168 17406
rect 284116 17342 284168 17348
rect 284680 10402 284708 84166
rect 284668 10396 284720 10402
rect 284668 10338 284720 10344
rect 283656 9036 283708 9042
rect 283656 8978 283708 8984
rect 284956 6322 284984 97854
rect 285140 84194 285168 100028
rect 285324 84194 285352 100028
rect 285508 84194 285536 100028
rect 285692 97510 285720 100028
rect 285680 97504 285732 97510
rect 285680 97446 285732 97452
rect 285876 96762 285904 100028
rect 286060 97306 286088 100028
rect 286048 97300 286100 97306
rect 286048 97242 286100 97248
rect 285864 96756 285916 96762
rect 285864 96698 285916 96704
rect 286244 84194 286272 100028
rect 286324 97980 286376 97986
rect 286324 97922 286376 97928
rect 285048 84166 285168 84194
rect 285232 84166 285352 84194
rect 285416 84166 285536 84194
rect 286152 84166 286272 84194
rect 285048 7682 285076 84166
rect 285232 7750 285260 84166
rect 285220 7744 285272 7750
rect 285220 7686 285272 7692
rect 285036 7676 285088 7682
rect 285036 7618 285088 7624
rect 284944 6316 284996 6322
rect 284944 6258 284996 6264
rect 285416 6186 285444 84166
rect 286152 10334 286180 84166
rect 286336 11762 286364 97922
rect 286324 11756 286376 11762
rect 286324 11698 286376 11704
rect 286140 10328 286192 10334
rect 286140 10270 286192 10276
rect 286428 6254 286456 100028
rect 286612 96898 286640 100028
rect 286600 96892 286652 96898
rect 286600 96834 286652 96840
rect 286796 84194 286824 100028
rect 286980 84194 287008 100028
rect 287164 97918 287192 100028
rect 287348 97986 287376 100028
rect 287336 97980 287388 97986
rect 287336 97922 287388 97928
rect 287152 97912 287204 97918
rect 287152 97854 287204 97860
rect 287152 96960 287204 96966
rect 287152 96902 287204 96908
rect 286704 84166 286824 84194
rect 286888 84166 287008 84194
rect 286704 9110 286732 84166
rect 286692 9104 286744 9110
rect 286692 9046 286744 9052
rect 286888 8974 286916 84166
rect 286876 8968 286928 8974
rect 286876 8910 286928 8916
rect 287164 7614 287192 96902
rect 287152 7608 287204 7614
rect 287152 7550 287204 7556
rect 286416 6248 286468 6254
rect 286416 6190 286468 6196
rect 285404 6180 285456 6186
rect 285404 6122 285456 6128
rect 285864 6180 285916 6186
rect 285864 6122 285916 6128
rect 283564 4956 283616 4962
rect 283564 4898 283616 4904
rect 282184 4888 282236 4894
rect 282184 4830 282236 4836
rect 282552 4480 282604 4486
rect 282552 4422 282604 4428
rect 281448 3800 281500 3806
rect 281448 3742 281500 3748
rect 281460 480 281488 3742
rect 282564 480 282592 4422
rect 284760 4004 284812 4010
rect 284760 3946 284812 3952
rect 283656 3868 283708 3874
rect 283656 3810 283708 3816
rect 283668 480 283696 3810
rect 284772 480 284800 3946
rect 285876 480 285904 6122
rect 286968 3936 287020 3942
rect 286968 3878 287020 3884
rect 286980 480 287008 3878
rect 287532 3466 287560 100028
rect 287716 96966 287744 100028
rect 287704 96960 287756 96966
rect 287704 96902 287756 96908
rect 287704 96756 287756 96762
rect 287704 96698 287756 96704
rect 287716 4486 287744 96698
rect 287900 84194 287928 100028
rect 288084 84194 288112 100028
rect 288268 84194 288296 100028
rect 288452 97442 288480 100028
rect 288440 97436 288492 97442
rect 288440 97378 288492 97384
rect 288636 96914 288664 100028
rect 288820 97850 288848 100028
rect 288808 97844 288860 97850
rect 288808 97786 288860 97792
rect 288636 96886 288940 96914
rect 288624 96824 288676 96830
rect 288624 96766 288676 96772
rect 287808 84166 287928 84194
rect 287992 84166 288112 84194
rect 288176 84166 288296 84194
rect 287808 63034 287836 84166
rect 287796 63028 287848 63034
rect 287796 62970 287848 62976
rect 287704 4480 287756 4486
rect 287704 4422 287756 4428
rect 287992 3534 288020 84166
rect 288176 5098 288204 84166
rect 288164 5092 288216 5098
rect 288164 5034 288216 5040
rect 288636 3670 288664 96766
rect 288624 3664 288676 3670
rect 288624 3606 288676 3612
rect 288912 3602 288940 96886
rect 289004 71058 289032 100028
rect 289188 97050 289216 100028
rect 289372 97578 289400 100028
rect 289360 97572 289412 97578
rect 289360 97514 289412 97520
rect 289096 97022 289216 97050
rect 289096 96830 289124 97022
rect 289176 96960 289228 96966
rect 289176 96902 289228 96908
rect 289084 96824 289136 96830
rect 289084 96766 289136 96772
rect 289084 96688 289136 96694
rect 289084 96630 289136 96636
rect 288992 71052 289044 71058
rect 288992 70994 289044 71000
rect 289096 5574 289124 96630
rect 289188 9178 289216 96902
rect 289556 84194 289584 100028
rect 289740 84194 289768 100028
rect 289924 96966 289952 100028
rect 289912 96960 289964 96966
rect 289912 96902 289964 96908
rect 290108 96694 290136 100028
rect 290096 96688 290148 96694
rect 290096 96630 290148 96636
rect 290292 84194 290320 100028
rect 290476 96762 290504 100028
rect 290464 96756 290516 96762
rect 290464 96698 290516 96704
rect 290660 84194 290688 100028
rect 290844 84194 290872 100028
rect 291028 84194 291056 100028
rect 291212 93854 291240 100028
rect 291396 96914 291424 100028
rect 291396 96886 291516 96914
rect 291212 93826 291424 93854
rect 289464 84166 289584 84194
rect 289648 84166 289768 84194
rect 290200 84166 290320 84194
rect 290568 84166 290688 84194
rect 290752 84166 290872 84194
rect 290936 84166 291056 84194
rect 289464 73846 289492 84166
rect 289452 73840 289504 73846
rect 289452 73782 289504 73788
rect 289176 9172 289228 9178
rect 289176 9114 289228 9120
rect 289084 5568 289136 5574
rect 289084 5510 289136 5516
rect 289648 3738 289676 84166
rect 290200 3806 290228 84166
rect 290568 3874 290596 84166
rect 290752 4010 290780 84166
rect 290936 6186 290964 84166
rect 290924 6180 290976 6186
rect 290924 6122 290976 6128
rect 290740 4004 290792 4010
rect 290740 3946 290792 3952
rect 291396 3942 291424 93826
rect 291384 3936 291436 3942
rect 291384 3878 291436 3884
rect 290556 3868 290608 3874
rect 290556 3810 290608 3816
rect 290188 3800 290240 3806
rect 290188 3742 290240 3748
rect 289636 3732 289688 3738
rect 289636 3674 289688 3680
rect 288900 3596 288952 3602
rect 288900 3538 288952 3544
rect 291488 3534 291516 96886
rect 287980 3528 288032 3534
rect 287980 3470 288032 3476
rect 288072 3528 288124 3534
rect 288072 3470 288124 3476
rect 291476 3528 291528 3534
rect 291476 3470 291528 3476
rect 287520 3460 287572 3466
rect 287520 3402 287572 3408
rect 288084 480 288112 3470
rect 290280 3460 290332 3466
rect 290280 3402 290332 3408
rect 289176 3188 289228 3194
rect 289176 3130 289228 3136
rect 289188 480 289216 3130
rect 290292 480 290320 3402
rect 291580 3194 291608 100028
rect 291764 3466 291792 100028
rect 291948 84194 291976 100028
rect 292132 84194 292160 100028
rect 292316 84194 292344 100028
rect 292500 84194 292528 100028
rect 292684 84194 292712 100028
rect 292868 84194 292896 100028
rect 293052 84194 293080 100028
rect 293236 84194 293264 100028
rect 293420 84194 293448 100028
rect 293604 84194 293632 100028
rect 293788 84194 293816 100028
rect 293972 97714 294000 100028
rect 294156 97850 294184 100028
rect 294144 97844 294196 97850
rect 294144 97786 294196 97792
rect 293960 97708 294012 97714
rect 293960 97650 294012 97656
rect 294340 97578 294368 100028
rect 294328 97572 294380 97578
rect 294328 97514 294380 97520
rect 294524 84194 294552 100028
rect 294708 84194 294736 100028
rect 294892 97782 294920 100028
rect 294880 97776 294932 97782
rect 294880 97718 294932 97724
rect 295076 84194 295104 100028
rect 295260 84194 295288 100028
rect 295444 84194 295472 100028
rect 295628 97646 295656 100028
rect 295616 97640 295668 97646
rect 295616 97582 295668 97588
rect 295812 84194 295840 100028
rect 295996 84194 296024 100028
rect 296180 84194 296208 100028
rect 296364 84194 296392 100028
rect 296548 84194 296576 100028
rect 291856 84166 291976 84194
rect 292040 84166 292160 84194
rect 292224 84166 292344 84194
rect 292408 84166 292528 84194
rect 292592 84166 292712 84194
rect 292776 84166 292896 84194
rect 292960 84166 293080 84194
rect 293144 84166 293264 84194
rect 293328 84166 293448 84194
rect 293512 84166 293632 84194
rect 293696 84166 293816 84194
rect 294432 84166 294552 84194
rect 294616 84166 294736 84194
rect 294984 84166 295104 84194
rect 295168 84166 295288 84194
rect 295352 84166 295472 84194
rect 295720 84166 295840 84194
rect 295904 84166 296024 84194
rect 296088 84166 296208 84194
rect 296272 84166 296392 84194
rect 296456 84166 296576 84194
rect 291752 3460 291804 3466
rect 291752 3402 291804 3408
rect 291568 3188 291620 3194
rect 291568 3130 291620 3136
rect 19770 -960 19882 480
rect 20874 -960 20986 480
rect 21978 -960 22090 480
rect 23082 -960 23194 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26394 -960 26506 480
rect 27498 -960 27610 480
rect 28602 -960 28714 480
rect 29706 -960 29818 480
rect 30810 -960 30922 480
rect 31914 -960 32026 480
rect 33018 -960 33130 480
rect 34122 -960 34234 480
rect 35226 -960 35338 480
rect 36330 -960 36442 480
rect 37434 -960 37546 480
rect 38538 -960 38650 480
rect 39642 -960 39754 480
rect 40746 -960 40858 480
rect 41850 -960 41962 480
rect 42954 -960 43066 480
rect 44058 -960 44170 480
rect 45162 -960 45274 480
rect 46266 -960 46378 480
rect 47370 -960 47482 480
rect 48474 -960 48586 480
rect 49578 -960 49690 480
rect 50682 -960 50794 480
rect 51786 -960 51898 480
rect 52890 -960 53002 480
rect 53994 -960 54106 480
rect 55098 -960 55210 480
rect 56202 -960 56314 480
rect 57306 -960 57418 480
rect 58410 -960 58522 480
rect 59514 -960 59626 480
rect 60618 -960 60730 480
rect 61722 -960 61834 480
rect 62826 -960 62938 480
rect 63930 -960 64042 480
rect 65034 -960 65146 480
rect 66138 -960 66250 480
rect 67242 -960 67354 480
rect 68346 -960 68458 480
rect 69450 -960 69562 480
rect 70554 -960 70666 480
rect 71658 -960 71770 480
rect 72762 -960 72874 480
rect 73866 -960 73978 480
rect 74970 -960 75082 480
rect 76074 -960 76186 480
rect 77178 -960 77290 480
rect 78282 -960 78394 480
rect 79386 -960 79498 480
rect 80490 -960 80602 480
rect 81594 -960 81706 480
rect 82698 -960 82810 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86010 -960 86122 480
rect 87114 -960 87226 480
rect 88218 -960 88330 480
rect 89322 -960 89434 480
rect 90426 -960 90538 480
rect 91530 -960 91642 480
rect 92634 -960 92746 480
rect 93738 -960 93850 480
rect 94842 -960 94954 480
rect 95946 -960 96058 480
rect 97050 -960 97162 480
rect 98154 -960 98266 480
rect 99258 -960 99370 480
rect 100362 -960 100474 480
rect 101466 -960 101578 480
rect 102570 -960 102682 480
rect 103674 -960 103786 480
rect 104778 -960 104890 480
rect 105882 -960 105994 480
rect 106986 -960 107098 480
rect 108090 -960 108202 480
rect 109194 -960 109306 480
rect 110298 -960 110410 480
rect 111402 -960 111514 480
rect 112506 -960 112618 480
rect 113610 -960 113722 480
rect 114714 -960 114826 480
rect 115818 -960 115930 480
rect 116922 -960 117034 480
rect 118026 -960 118138 480
rect 119130 -960 119242 480
rect 120234 -960 120346 480
rect 121338 -960 121450 480
rect 122442 -960 122554 480
rect 123546 -960 123658 480
rect 124650 -960 124762 480
rect 125754 -960 125866 480
rect 126858 -960 126970 480
rect 127962 -960 128074 480
rect 129066 -960 129178 480
rect 130170 -960 130282 480
rect 131274 -960 131386 480
rect 132378 -960 132490 480
rect 133482 -960 133594 480
rect 134586 -960 134698 480
rect 135690 -960 135802 480
rect 136794 -960 136906 480
rect 137898 -960 138010 480
rect 139002 -960 139114 480
rect 140106 -960 140218 480
rect 141210 -960 141322 480
rect 142314 -960 142426 480
rect 143418 -960 143530 480
rect 144522 -960 144634 480
rect 145626 -960 145738 480
rect 146730 -960 146842 480
rect 147834 -960 147946 480
rect 148938 -960 149050 480
rect 150042 -960 150154 480
rect 151146 -960 151258 480
rect 152250 -960 152362 480
rect 153354 -960 153466 480
rect 154458 -960 154570 480
rect 155562 -960 155674 480
rect 156666 -960 156778 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 159978 -960 160090 480
rect 161082 -960 161194 480
rect 162186 -960 162298 480
rect 163290 -960 163402 480
rect 164394 -960 164506 480
rect 165498 -960 165610 480
rect 166602 -960 166714 480
rect 167706 -960 167818 480
rect 168810 -960 168922 480
rect 169914 -960 170026 480
rect 171018 -960 171130 480
rect 172122 -960 172234 480
rect 173226 -960 173338 480
rect 174330 -960 174442 480
rect 175434 -960 175546 480
rect 176538 -960 176650 480
rect 177642 -960 177754 480
rect 178746 -960 178858 480
rect 179850 -960 179962 480
rect 180954 -960 181066 480
rect 182058 -960 182170 480
rect 183162 -960 183274 480
rect 184266 -960 184378 480
rect 185370 -960 185482 480
rect 186474 -960 186586 480
rect 187578 -960 187690 480
rect 188682 -960 188794 480
rect 189786 -960 189898 480
rect 190890 -960 191002 480
rect 191994 -960 192106 480
rect 193098 -960 193210 480
rect 194202 -960 194314 480
rect 195306 -960 195418 480
rect 196410 -960 196522 480
rect 197514 -960 197626 480
rect 198618 -960 198730 480
rect 199722 -960 199834 480
rect 200826 -960 200938 480
rect 201930 -960 202042 480
rect 203034 -960 203146 480
rect 204138 -960 204250 480
rect 205242 -960 205354 480
rect 206346 -960 206458 480
rect 207450 -960 207562 480
rect 208554 -960 208666 480
rect 209658 -960 209770 480
rect 210762 -960 210874 480
rect 211866 -960 211978 480
rect 212970 -960 213082 480
rect 214074 -960 214186 480
rect 215178 -960 215290 480
rect 216282 -960 216394 480
rect 217386 -960 217498 480
rect 218490 -960 218602 480
rect 219594 -960 219706 480
rect 220698 -960 220810 480
rect 221802 -960 221914 480
rect 222906 -960 223018 480
rect 224010 -960 224122 480
rect 225114 -960 225226 480
rect 226218 -960 226330 480
rect 227322 -960 227434 480
rect 228426 -960 228538 480
rect 229530 -960 229642 480
rect 230634 -960 230746 480
rect 231738 -960 231850 480
rect 232842 -960 232954 480
rect 233946 -960 234058 480
rect 235050 -960 235162 480
rect 236154 -960 236266 480
rect 237258 -960 237370 480
rect 238362 -960 238474 480
rect 239466 -960 239578 480
rect 240570 -960 240682 480
rect 241674 -960 241786 480
rect 242778 -960 242890 480
rect 243882 -960 243994 480
rect 244986 -960 245098 480
rect 246090 -960 246202 480
rect 247194 -960 247306 480
rect 248298 -960 248410 480
rect 249402 -960 249514 480
rect 250506 -960 250618 480
rect 251610 -960 251722 480
rect 252714 -960 252826 480
rect 253818 -960 253930 480
rect 254922 -960 255034 480
rect 256026 -960 256138 480
rect 257130 -960 257242 480
rect 258234 -960 258346 480
rect 259338 -960 259450 480
rect 260442 -960 260554 480
rect 261546 -960 261658 480
rect 262650 -960 262762 480
rect 263754 -960 263866 480
rect 264858 -960 264970 480
rect 265962 -960 266074 480
rect 267066 -960 267178 480
rect 268170 -960 268282 480
rect 269274 -960 269386 480
rect 270378 -960 270490 480
rect 271482 -960 271594 480
rect 272586 -960 272698 480
rect 273690 -960 273802 480
rect 274794 -960 274906 480
rect 275898 -960 276010 480
rect 277002 -960 277114 480
rect 278106 -960 278218 480
rect 279210 -960 279322 480
rect 280314 -960 280426 480
rect 281418 -960 281530 480
rect 282522 -960 282634 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285834 -960 285946 480
rect 286938 -960 287050 480
rect 288042 -960 288154 480
rect 289146 -960 289258 480
rect 290250 -960 290362 480
rect 291354 354 291466 480
rect 291856 354 291884 84166
rect 292040 16574 292068 84166
rect 292040 16546 292160 16574
rect 292132 3482 292160 16546
rect 292224 3602 292252 84166
rect 292408 3670 292436 84166
rect 292396 3664 292448 3670
rect 292396 3606 292448 3612
rect 292212 3596 292264 3602
rect 292212 3538 292264 3544
rect 292132 3454 292528 3482
rect 292500 480 292528 3454
rect 292592 3398 292620 84166
rect 292776 3942 292804 84166
rect 292960 4146 292988 84166
rect 293144 4418 293172 84166
rect 293328 10334 293356 84166
rect 293316 10328 293368 10334
rect 293316 10270 293368 10276
rect 293132 4412 293184 4418
rect 293132 4354 293184 4360
rect 292948 4140 293000 4146
rect 292948 4082 293000 4088
rect 292764 3936 292816 3942
rect 292764 3878 292816 3884
rect 293512 3466 293540 84166
rect 293696 4962 293724 84166
rect 294432 83502 294460 84166
rect 294420 83496 294472 83502
rect 294420 83438 294472 83444
rect 294616 6254 294644 84166
rect 294984 69698 295012 84166
rect 294972 69692 295024 69698
rect 294972 69634 295024 69640
rect 295168 14482 295196 84166
rect 295156 14476 295208 14482
rect 295156 14418 295208 14424
rect 294604 6248 294656 6254
rect 294604 6190 294656 6196
rect 293684 4956 293736 4962
rect 293684 4898 293736 4904
rect 295352 4894 295380 84166
rect 295720 60042 295748 84166
rect 295708 60036 295760 60042
rect 295708 59978 295760 59984
rect 295904 6186 295932 84166
rect 295892 6180 295944 6186
rect 295892 6122 295944 6128
rect 295340 4888 295392 4894
rect 295340 4830 295392 4836
rect 296088 4826 296116 84166
rect 296272 62830 296300 84166
rect 296260 62824 296312 62830
rect 296260 62766 296312 62772
rect 296456 7614 296484 84166
rect 296732 9042 296760 100028
rect 296916 84194 296944 100028
rect 297100 97374 297128 100028
rect 297088 97368 297140 97374
rect 297088 97310 297140 97316
rect 297284 84194 297312 100028
rect 297468 84194 297496 100028
rect 297652 97306 297680 100028
rect 297640 97300 297692 97306
rect 297640 97242 297692 97248
rect 297836 84194 297864 100028
rect 298020 84194 298048 100028
rect 298204 97442 298232 100028
rect 298192 97436 298244 97442
rect 298192 97378 298244 97384
rect 298388 84194 298416 100028
rect 298572 84194 298600 100028
rect 298756 94518 298784 100028
rect 298744 94512 298796 94518
rect 298744 94454 298796 94460
rect 298940 84194 298968 100028
rect 299124 84194 299152 100028
rect 299308 97510 299336 100028
rect 299296 97504 299348 97510
rect 299296 97446 299348 97452
rect 296824 84166 296944 84194
rect 297192 84166 297312 84194
rect 297376 84166 297496 84194
rect 297744 84166 297864 84194
rect 297928 84166 298048 84194
rect 298296 84166 298416 84194
rect 298480 84166 298600 84194
rect 298848 84166 298968 84194
rect 299032 84166 299152 84194
rect 296824 64190 296852 84166
rect 296812 64184 296864 64190
rect 296812 64126 296864 64132
rect 297192 54534 297220 84166
rect 297180 54528 297232 54534
rect 297180 54470 297232 54476
rect 297376 32434 297404 84166
rect 297364 32428 297416 32434
rect 297364 32370 297416 32376
rect 297744 11762 297772 84166
rect 297928 44878 297956 84166
rect 297916 44872 297968 44878
rect 297916 44814 297968 44820
rect 298296 13122 298324 84166
rect 298480 46238 298508 84166
rect 298848 72486 298876 84166
rect 298836 72480 298888 72486
rect 298836 72422 298888 72428
rect 298468 46232 298520 46238
rect 298468 46174 298520 46180
rect 299032 35290 299060 84166
rect 299492 61538 299520 100028
rect 299676 84194 299704 100028
rect 299860 96286 299888 100028
rect 299848 96280 299900 96286
rect 299848 96222 299900 96228
rect 300044 90642 300072 100028
rect 300228 96914 300256 100028
rect 300308 97844 300360 97850
rect 300308 97786 300360 97792
rect 300136 96886 300256 96914
rect 300032 90636 300084 90642
rect 300032 90578 300084 90584
rect 299584 84166 299704 84194
rect 299480 61532 299532 61538
rect 299480 61474 299532 61480
rect 299020 35284 299072 35290
rect 299020 35226 299072 35232
rect 299584 22846 299612 84166
rect 300136 80918 300164 96886
rect 300320 96778 300348 97786
rect 300228 96750 300348 96778
rect 300124 80912 300176 80918
rect 300124 80854 300176 80860
rect 299572 22840 299624 22846
rect 299572 22782 299624 22788
rect 298284 13116 298336 13122
rect 298284 13058 298336 13064
rect 297732 11756 297784 11762
rect 297732 11698 297784 11704
rect 300228 11014 300256 96750
rect 300412 91934 300440 100028
rect 300400 91928 300452 91934
rect 300400 91870 300452 91876
rect 300596 84194 300624 100028
rect 300780 84194 300808 100028
rect 300860 97708 300912 97714
rect 300860 97650 300912 97656
rect 300872 96762 300900 97650
rect 300860 96756 300912 96762
rect 300860 96698 300912 96704
rect 300964 93362 300992 100028
rect 301148 96830 301176 100028
rect 301136 96824 301188 96830
rect 301136 96766 301188 96772
rect 300952 93356 301004 93362
rect 300952 93298 301004 93304
rect 301332 84194 301360 100028
rect 301516 96914 301544 100028
rect 301700 96914 301728 100028
rect 301780 97776 301832 97782
rect 301780 97718 301832 97724
rect 301424 96886 301544 96914
rect 301608 96886 301728 96914
rect 301424 89282 301452 96886
rect 301504 96756 301556 96762
rect 301504 96698 301556 96704
rect 301412 89276 301464 89282
rect 301412 89218 301464 89224
rect 300504 84166 300624 84194
rect 300688 84166 300808 84194
rect 301240 84166 301360 84194
rect 300504 76770 300532 84166
rect 300492 76764 300544 76770
rect 300492 76706 300544 76712
rect 300216 11008 300268 11014
rect 300216 10950 300268 10956
rect 300688 10334 300716 84166
rect 301240 40866 301268 84166
rect 301228 40860 301280 40866
rect 301228 40802 301280 40808
rect 300216 10328 300268 10334
rect 300216 10270 300268 10276
rect 300676 10328 300728 10334
rect 300676 10270 300728 10276
rect 296720 9036 296772 9042
rect 296720 8978 296772 8984
rect 296444 7608 296496 7614
rect 296444 7550 296496 7556
rect 296076 4820 296128 4826
rect 296076 4762 296128 4768
rect 299112 4412 299164 4418
rect 299112 4354 299164 4360
rect 298008 4140 298060 4146
rect 298008 4082 298060 4088
rect 296904 3936 296956 3942
rect 296904 3878 296956 3884
rect 294696 3664 294748 3670
rect 294696 3606 294748 3612
rect 293592 3596 293644 3602
rect 293592 3538 293644 3544
rect 293500 3460 293552 3466
rect 293500 3402 293552 3408
rect 292580 3392 292632 3398
rect 292580 3334 292632 3340
rect 293604 480 293632 3538
rect 294708 480 294736 3606
rect 295800 3392 295852 3398
rect 295800 3334 295852 3340
rect 295812 480 295840 3334
rect 296916 480 296944 3878
rect 298020 480 298048 4082
rect 299124 480 299152 4354
rect 300228 480 300256 10270
rect 301516 4214 301544 96698
rect 301608 75342 301636 96886
rect 301792 96778 301820 97718
rect 301700 96750 301820 96778
rect 301596 75336 301648 75342
rect 301596 75278 301648 75284
rect 301700 4554 301728 96750
rect 301884 84194 301912 100028
rect 302068 87854 302096 100028
rect 302056 87848 302108 87854
rect 302056 87790 302108 87796
rect 301792 84166 301912 84194
rect 301792 82346 301820 84166
rect 301780 82340 301832 82346
rect 301780 82282 301832 82288
rect 302252 79558 302280 100028
rect 302436 84194 302464 100028
rect 302620 96218 302648 100028
rect 302608 96212 302660 96218
rect 302608 96154 302660 96160
rect 302804 84194 302832 100028
rect 302988 96914 303016 100028
rect 302344 84166 302464 84194
rect 302712 84166 302832 84194
rect 302896 96886 303016 96914
rect 302240 79552 302292 79558
rect 302240 79494 302292 79500
rect 302344 33930 302372 84166
rect 302712 72690 302740 84166
rect 302700 72684 302752 72690
rect 302700 72626 302752 72632
rect 302332 33924 302384 33930
rect 302332 33866 302384 33872
rect 302896 8974 302924 96886
rect 302976 96824 303028 96830
rect 302976 96766 303028 96772
rect 302988 93430 303016 96766
rect 303172 94790 303200 100028
rect 303160 94784 303212 94790
rect 303160 94726 303212 94732
rect 302976 93424 303028 93430
rect 302976 93366 303028 93372
rect 303356 84194 303384 100028
rect 303540 84194 303568 100028
rect 303620 97572 303672 97578
rect 303620 97514 303672 97520
rect 303632 96830 303660 97514
rect 303620 96824 303672 96830
rect 303620 96766 303672 96772
rect 303724 92070 303752 100028
rect 303908 97986 303936 100028
rect 303896 97980 303948 97986
rect 303896 97922 303948 97928
rect 303712 92064 303764 92070
rect 303712 92006 303764 92012
rect 304092 84194 304120 100028
rect 304276 96914 304304 100028
rect 304460 96914 304488 100028
rect 304540 97640 304592 97646
rect 304540 97582 304592 97588
rect 304184 96886 304304 96914
rect 304368 96886 304488 96914
rect 304184 90506 304212 96886
rect 304264 96824 304316 96830
rect 304264 96766 304316 96772
rect 304172 90500 304224 90506
rect 304172 90442 304224 90448
rect 303264 84166 303384 84194
rect 303448 84166 303568 84194
rect 304000 84166 304120 84194
rect 303264 78198 303292 84166
rect 303252 78192 303304 78198
rect 303252 78134 303304 78140
rect 303448 39506 303476 84166
rect 304000 67046 304028 84166
rect 303988 67040 304040 67046
rect 303988 66982 304040 66988
rect 303436 39500 303488 39506
rect 303436 39442 303488 39448
rect 304172 11008 304224 11014
rect 304172 10950 304224 10956
rect 302884 8968 302936 8974
rect 302884 8910 302936 8916
rect 302424 4956 302476 4962
rect 302424 4898 302476 4904
rect 301688 4548 301740 4554
rect 301688 4490 301740 4496
rect 301504 4208 301556 4214
rect 301504 4150 301556 4156
rect 301320 3460 301372 3466
rect 301320 3402 301372 3408
rect 301332 480 301360 3402
rect 302436 480 302464 4898
rect 303528 4208 303580 4214
rect 303528 4150 303580 4156
rect 303540 480 303568 4150
rect 304184 3482 304212 10950
rect 304276 4214 304304 96766
rect 304368 61470 304396 96886
rect 304552 96778 304580 97582
rect 304460 96750 304580 96778
rect 304356 61464 304408 61470
rect 304356 61406 304408 61412
rect 304460 6322 304488 96750
rect 304644 84194 304672 100028
rect 304828 86494 304856 100028
rect 304816 86488 304868 86494
rect 304816 86430 304868 86436
rect 304552 84166 304672 84194
rect 304552 38010 304580 84166
rect 305012 73982 305040 100028
rect 305196 84194 305224 100028
rect 305380 89214 305408 100028
rect 305368 89208 305420 89214
rect 305368 89150 305420 89156
rect 305564 84194 305592 100028
rect 305748 84194 305776 100028
rect 305932 87786 305960 100028
rect 305920 87780 305972 87786
rect 305920 87722 305972 87728
rect 306116 84194 306144 100028
rect 306300 84194 306328 100028
rect 306484 85066 306512 100028
rect 306472 85060 306524 85066
rect 306472 85002 306524 85008
rect 306668 84194 306696 100028
rect 306852 84194 306880 100028
rect 307036 96914 307064 100028
rect 307116 97980 307168 97986
rect 307116 97922 307168 97928
rect 305104 84166 305224 84194
rect 305472 84166 305592 84194
rect 305656 84166 305776 84194
rect 306024 84166 306144 84194
rect 306208 84166 306328 84194
rect 306576 84166 306696 84194
rect 306760 84166 306880 84194
rect 306944 96886 307064 96914
rect 305000 73976 305052 73982
rect 305000 73918 305052 73924
rect 304540 38004 304592 38010
rect 304540 37946 304592 37952
rect 305104 36650 305132 84166
rect 305472 76702 305500 84166
rect 305460 76696 305512 76702
rect 305460 76638 305512 76644
rect 305092 36644 305144 36650
rect 305092 36586 305144 36592
rect 305656 7682 305684 84166
rect 306024 49094 306052 84166
rect 306012 49088 306064 49094
rect 306012 49030 306064 49036
rect 306208 35222 306236 84166
rect 306380 83496 306432 83502
rect 306380 83438 306432 83444
rect 306196 35216 306248 35222
rect 306196 35158 306248 35164
rect 305644 7676 305696 7682
rect 305644 7618 305696 7624
rect 306392 6914 306420 83438
rect 306576 58818 306604 84166
rect 306564 58812 306616 58818
rect 306564 58754 306616 58760
rect 306760 11830 306788 84166
rect 306944 83706 306972 96886
rect 307128 96778 307156 97922
rect 307036 96750 307156 96778
rect 307036 90574 307064 96750
rect 307024 90568 307076 90574
rect 307024 90510 307076 90516
rect 307220 84194 307248 100028
rect 307404 84194 307432 100028
rect 307588 84194 307616 100028
rect 307772 86426 307800 100028
rect 307956 92002 307984 100028
rect 308140 96830 308168 100028
rect 308128 96824 308180 96830
rect 308128 96766 308180 96772
rect 307944 91996 307996 92002
rect 307944 91938 307996 91944
rect 308324 87718 308352 100028
rect 308312 87712 308364 87718
rect 308312 87654 308364 87660
rect 307760 86420 307812 86426
rect 307760 86362 307812 86368
rect 308508 84194 308536 100028
rect 308692 96150 308720 100028
rect 308680 96144 308732 96150
rect 308680 96086 308732 96092
rect 308876 84194 308904 100028
rect 309060 84194 309088 100028
rect 309244 84194 309272 100028
rect 309428 84194 309456 100028
rect 309612 84194 309640 100028
rect 309796 96914 309824 100028
rect 307128 84166 307248 84194
rect 307312 84166 307432 84194
rect 307496 84166 307616 84194
rect 308416 84166 308536 84194
rect 308784 84166 308904 84194
rect 308968 84166 309088 84194
rect 309152 84166 309272 84194
rect 309336 84166 309456 84194
rect 309520 84166 309640 84194
rect 309704 96886 309824 96914
rect 306932 83700 306984 83706
rect 306932 83642 306984 83648
rect 307128 57390 307156 84166
rect 307116 57384 307168 57390
rect 307116 57326 307168 57332
rect 307312 22778 307340 84166
rect 307496 80850 307524 84166
rect 307484 80844 307536 80850
rect 307484 80786 307536 80792
rect 308416 32502 308444 84166
rect 308784 72622 308812 84166
rect 308772 72616 308824 72622
rect 308772 72558 308824 72564
rect 308404 32496 308456 32502
rect 308404 32438 308456 32444
rect 307300 22772 307352 22778
rect 307300 22714 307352 22720
rect 308968 13190 308996 84166
rect 309152 82278 309180 84166
rect 309140 82272 309192 82278
rect 309140 82214 309192 82220
rect 309140 69692 309192 69698
rect 309140 69634 309192 69640
rect 308956 13184 309008 13190
rect 308956 13126 309008 13132
rect 306748 11824 306800 11830
rect 306748 11766 306800 11772
rect 309152 6914 309180 69634
rect 309336 56030 309364 84166
rect 309520 65686 309548 84166
rect 309704 71194 309732 96886
rect 309784 96824 309836 96830
rect 309784 96766 309836 96772
rect 309796 93294 309824 96766
rect 309784 93288 309836 93294
rect 309784 93230 309836 93236
rect 309980 84194 310008 100028
rect 310164 84194 310192 100028
rect 310348 84194 310376 100028
rect 309888 84166 310008 84194
rect 310072 84166 310192 84194
rect 310256 84166 310376 84194
rect 309692 71188 309744 71194
rect 309692 71130 309744 71136
rect 309508 65680 309560 65686
rect 309508 65622 309560 65628
rect 309324 56024 309376 56030
rect 309324 55966 309376 55972
rect 309888 51814 309916 84166
rect 309876 51808 309928 51814
rect 309876 51750 309928 51756
rect 310072 10402 310100 84166
rect 310256 69834 310284 84166
rect 310244 69828 310296 69834
rect 310244 69770 310296 69776
rect 310532 53174 310560 100028
rect 310716 94722 310744 100028
rect 310704 94716 310756 94722
rect 310704 94658 310756 94664
rect 310900 86358 310928 100028
rect 310888 86352 310940 86358
rect 310888 86294 310940 86300
rect 311084 84194 311112 100028
rect 311268 84194 311296 100028
rect 311452 84194 311480 100028
rect 311636 84194 311664 100028
rect 311820 84194 311848 100028
rect 312004 96830 312032 100028
rect 311992 96824 312044 96830
rect 311992 96766 312044 96772
rect 312188 84998 312216 100028
rect 312176 84992 312228 84998
rect 312176 84934 312228 84940
rect 312372 84194 312400 100028
rect 312556 87650 312584 100028
rect 312544 87644 312596 87650
rect 312544 87586 312596 87592
rect 312740 84194 312768 100028
rect 312924 84194 312952 100028
rect 313108 84194 313136 100028
rect 310992 84166 311112 84194
rect 311176 84166 311296 84194
rect 311360 84166 311480 84194
rect 311544 84166 311664 84194
rect 311728 84166 311848 84194
rect 312280 84166 312400 84194
rect 312648 84166 312768 84194
rect 312832 84166 312952 84194
rect 313016 84166 313136 84194
rect 310992 75274 311020 84166
rect 310980 75268 311032 75274
rect 310980 75210 311032 75216
rect 310520 53168 310572 53174
rect 310520 53110 310572 53116
rect 311176 40798 311204 84166
rect 311360 79490 311388 84166
rect 311348 79484 311400 79490
rect 311348 79426 311400 79432
rect 311164 40792 311216 40798
rect 311164 40734 311216 40740
rect 311544 31142 311572 84166
rect 311728 49026 311756 84166
rect 312280 62966 312308 84166
rect 312268 62960 312320 62966
rect 312268 62902 312320 62908
rect 311716 49020 311768 49026
rect 311716 48962 311768 48968
rect 311532 31136 311584 31142
rect 311532 31078 311584 31084
rect 312648 29714 312676 84166
rect 312832 39438 312860 84166
rect 313016 78130 313044 84166
rect 313292 79422 313320 100028
rect 313476 84194 313504 100028
rect 313660 94654 313688 100028
rect 313648 94648 313700 94654
rect 313648 94590 313700 94596
rect 313844 84194 313872 100028
rect 314028 84194 314056 100028
rect 314212 84194 314240 100028
rect 314396 84194 314424 100028
rect 314580 84194 314608 100028
rect 314764 84930 314792 100028
rect 314752 84924 314804 84930
rect 314752 84866 314804 84872
rect 314948 84194 314976 100028
rect 315132 84194 315160 100028
rect 315316 96914 315344 100028
rect 313384 84166 313504 84194
rect 313752 84166 313872 84194
rect 313936 84166 314056 84194
rect 314120 84166 314240 84194
rect 314304 84166 314424 84194
rect 314488 84166 314608 84194
rect 314856 84166 314976 84194
rect 315040 84166 315160 84194
rect 315224 96886 315344 96914
rect 313280 79416 313332 79422
rect 313280 79358 313332 79364
rect 313004 78124 313056 78130
rect 313004 78066 313056 78072
rect 313384 60178 313412 84166
rect 313372 60172 313424 60178
rect 313372 60114 313424 60120
rect 313280 60036 313332 60042
rect 313280 59978 313332 59984
rect 312820 39432 312872 39438
rect 312820 39374 312872 39380
rect 312636 29708 312688 29714
rect 312636 29650 312688 29656
rect 311256 14476 311308 14482
rect 311256 14418 311308 14424
rect 310060 10396 310112 10402
rect 310060 10338 310112 10344
rect 306392 6886 306880 6914
rect 309152 6886 310192 6914
rect 304448 6316 304500 6322
rect 304448 6258 304500 6264
rect 304264 4208 304316 4214
rect 304264 4150 304316 4156
rect 305736 4208 305788 4214
rect 305736 4150 305788 4156
rect 304184 3454 304672 3482
rect 304644 480 304672 3454
rect 305748 480 305776 4150
rect 306852 480 306880 6886
rect 307944 6248 307996 6254
rect 307944 6190 307996 6196
rect 307956 480 307984 6190
rect 309048 4548 309100 4554
rect 309048 4490 309100 4496
rect 309060 480 309088 4490
rect 310164 480 310192 6886
rect 311268 480 311296 14418
rect 312360 4888 312412 4894
rect 312360 4830 312412 4836
rect 312372 480 312400 4830
rect 313292 3534 313320 59978
rect 313752 54602 313780 84166
rect 313740 54596 313792 54602
rect 313740 54538 313792 54544
rect 313936 33862 313964 84166
rect 314120 75206 314148 84166
rect 314108 75200 314160 75206
rect 314108 75142 314160 75148
rect 313924 33856 313976 33862
rect 313924 33798 313976 33804
rect 314304 28354 314332 84166
rect 314488 64326 314516 84166
rect 314476 64320 314528 64326
rect 314476 64262 314528 64268
rect 314292 28348 314344 28354
rect 314292 28290 314344 28296
rect 314856 26994 314884 84166
rect 314844 26988 314896 26994
rect 314844 26930 314896 26936
rect 313464 6316 313516 6322
rect 313464 6258 313516 6264
rect 313280 3528 313332 3534
rect 313280 3470 313332 3476
rect 313476 480 313504 6258
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 314580 480 314608 3470
rect 315040 3262 315068 84166
rect 315224 68474 315252 96886
rect 315304 96824 315356 96830
rect 315304 96766 315356 96772
rect 315316 89146 315344 96766
rect 315304 89140 315356 89146
rect 315304 89082 315356 89088
rect 315500 84194 315528 100028
rect 315684 84194 315712 100028
rect 315868 84194 315896 100028
rect 316052 96082 316080 100028
rect 316040 96076 316092 96082
rect 316040 96018 316092 96024
rect 316236 84194 316264 100028
rect 316420 97714 316448 100028
rect 316408 97708 316460 97714
rect 316408 97650 316460 97656
rect 316604 84194 316632 100028
rect 316788 84194 316816 100028
rect 316972 96830 317000 100028
rect 316960 96824 317012 96830
rect 316960 96766 317012 96772
rect 317156 84194 317184 100028
rect 317340 84194 317368 100028
rect 317524 84194 317552 100028
rect 317708 84194 317736 100028
rect 317892 84194 317920 100028
rect 318076 96914 318104 100028
rect 315408 84166 315528 84194
rect 315592 84166 315712 84194
rect 315776 84166 315896 84194
rect 316144 84166 316264 84194
rect 316512 84166 316632 84194
rect 316696 84166 316816 84194
rect 317064 84166 317184 84194
rect 317248 84166 317368 84194
rect 317432 84166 317552 84194
rect 317616 84166 317736 84194
rect 317800 84166 317920 84194
rect 317984 96886 318104 96914
rect 315212 68468 315264 68474
rect 315212 68410 315264 68416
rect 315408 25634 315436 84166
rect 315396 25628 315448 25634
rect 315396 25570 315448 25576
rect 315592 3330 315620 84166
rect 315776 66978 315804 84166
rect 315764 66972 315816 66978
rect 315764 66914 315816 66920
rect 315672 6180 315724 6186
rect 315672 6122 315724 6128
rect 315580 3324 315632 3330
rect 315580 3266 315632 3272
rect 315028 3256 315080 3262
rect 315028 3198 315080 3204
rect 315684 480 315712 6122
rect 316144 3398 316172 84166
rect 316512 71126 316540 84166
rect 316500 71120 316552 71126
rect 316500 71062 316552 71068
rect 316696 4146 316724 84166
rect 317064 78062 317092 84166
rect 317052 78056 317104 78062
rect 317052 77998 317104 78004
rect 316776 4820 316828 4826
rect 316776 4762 316828 4768
rect 316684 4140 316736 4146
rect 316684 4082 316736 4088
rect 316132 3392 316184 3398
rect 316132 3334 316184 3340
rect 316788 480 316816 4762
rect 317248 4078 317276 84166
rect 317432 65618 317460 84166
rect 317420 65612 317472 65618
rect 317420 65554 317472 65560
rect 317420 62824 317472 62830
rect 317420 62766 317472 62772
rect 317432 16574 317460 62766
rect 317616 24206 317644 84166
rect 317604 24200 317656 24206
rect 317604 24142 317656 24148
rect 317432 16546 317736 16574
rect 317236 4072 317288 4078
rect 317236 4014 317288 4020
rect 317708 3482 317736 16546
rect 317800 4010 317828 84166
rect 317984 64258 318012 96886
rect 318064 96824 318116 96830
rect 318064 96766 318116 96772
rect 318076 83638 318104 96766
rect 318260 84194 318288 100028
rect 318444 84194 318472 100028
rect 318628 84194 318656 100028
rect 318812 96762 318840 100028
rect 318800 96756 318852 96762
rect 318800 96698 318852 96704
rect 318996 84194 319024 100028
rect 319180 91866 319208 100028
rect 319168 91860 319220 91866
rect 319168 91802 319220 91808
rect 319364 84194 319392 100028
rect 319548 84194 319576 100028
rect 319732 84194 319760 100028
rect 319916 84194 319944 100028
rect 320100 84194 320128 100028
rect 320284 84194 320312 100028
rect 320468 84194 320496 100028
rect 320652 84194 320680 100028
rect 320836 96914 320864 100028
rect 320916 97368 320968 97374
rect 320916 97310 320968 97316
rect 318168 84166 318288 84194
rect 318352 84166 318472 84194
rect 318536 84166 318656 84194
rect 318904 84166 319024 84194
rect 319272 84166 319392 84194
rect 319456 84166 319576 84194
rect 319640 84166 319760 84194
rect 319824 84166 319944 84194
rect 320008 84166 320128 84194
rect 320192 84166 320312 84194
rect 320376 84166 320496 84194
rect 320560 84166 320680 84194
rect 320744 96886 320864 96914
rect 318064 83632 318116 83638
rect 318064 83574 318116 83580
rect 317972 64252 318024 64258
rect 317972 64194 318024 64200
rect 318168 21486 318196 84166
rect 318156 21480 318208 21486
rect 318156 21422 318208 21428
rect 317788 4004 317840 4010
rect 317788 3946 317840 3952
rect 318352 3942 318380 84166
rect 318536 62898 318564 84166
rect 318524 62892 318576 62898
rect 318524 62834 318576 62840
rect 318340 3936 318392 3942
rect 318340 3878 318392 3884
rect 318904 3874 318932 84166
rect 319272 61402 319300 84166
rect 319260 61396 319312 61402
rect 319260 61338 319312 61344
rect 318984 7608 319036 7614
rect 318984 7550 319036 7556
rect 318892 3868 318944 3874
rect 318892 3810 318944 3816
rect 317708 3454 317920 3482
rect 317892 480 317920 3454
rect 318996 480 319024 7550
rect 319456 3806 319484 84166
rect 319640 71058 319668 84166
rect 319628 71052 319680 71058
rect 319628 70994 319680 71000
rect 319824 20058 319852 84166
rect 319812 20052 319864 20058
rect 319812 19994 319864 20000
rect 319444 3800 319496 3806
rect 319444 3742 319496 3748
rect 320008 3738 320036 84166
rect 320192 69766 320220 84166
rect 320376 83570 320404 84166
rect 320364 83564 320416 83570
rect 320364 83506 320416 83512
rect 320180 69760 320232 69766
rect 320180 69702 320232 69708
rect 320180 64184 320232 64190
rect 320180 64126 320232 64132
rect 320192 16574 320220 64126
rect 320192 16546 320496 16574
rect 320088 9036 320140 9042
rect 320088 8978 320140 8984
rect 319996 3732 320048 3738
rect 319996 3674 320048 3680
rect 320100 480 320128 8978
rect 320468 3482 320496 16546
rect 320560 3670 320588 84166
rect 320744 60110 320772 96886
rect 320928 96778 320956 97310
rect 320836 96750 320956 96778
rect 320732 60104 320784 60110
rect 320732 60046 320784 60052
rect 320836 4214 320864 96750
rect 321020 84194 321048 100028
rect 321204 84194 321232 100028
rect 321388 97374 321416 100028
rect 321376 97368 321428 97374
rect 321376 97310 321428 97316
rect 320928 84166 321048 84194
rect 321112 84166 321232 84194
rect 320928 18698 320956 84166
rect 320916 18692 320968 18698
rect 320916 18634 320968 18640
rect 321112 16574 321140 84166
rect 321572 73914 321600 100028
rect 321756 84194 321784 100028
rect 321940 97646 321968 100028
rect 321928 97640 321980 97646
rect 321928 97582 321980 97588
rect 322124 84194 322152 100028
rect 322308 84194 322336 100028
rect 322492 97578 322520 100028
rect 322480 97572 322532 97578
rect 322480 97514 322532 97520
rect 322676 84194 322704 100028
rect 322860 84194 322888 100028
rect 322940 97504 322992 97510
rect 322940 97446 322992 97452
rect 322952 96830 322980 97446
rect 322940 96824 322992 96830
rect 322940 96766 322992 96772
rect 323044 96014 323072 100028
rect 323032 96008 323084 96014
rect 323032 95950 323084 95956
rect 323228 84194 323256 100028
rect 323412 84194 323440 100028
rect 323492 97300 323544 97306
rect 323492 97242 323544 97248
rect 323504 93854 323532 97242
rect 323596 94586 323624 100028
rect 323780 96914 323808 100028
rect 323964 96914 323992 100028
rect 324044 97436 324096 97442
rect 324044 97378 324096 97384
rect 323688 96886 323808 96914
rect 323872 96886 323992 96914
rect 323584 94580 323636 94586
rect 323584 94522 323636 94528
rect 323504 93826 323624 93854
rect 321664 84166 321784 84194
rect 322032 84166 322152 84194
rect 322216 84166 322336 84194
rect 322584 84166 322704 84194
rect 322768 84166 322888 84194
rect 323136 84166 323256 84194
rect 323320 84166 323440 84194
rect 321560 73908 321612 73914
rect 321560 73850 321612 73856
rect 321664 17338 321692 84166
rect 322032 58750 322060 84166
rect 322020 58744 322072 58750
rect 322020 58686 322072 58692
rect 321652 17332 321704 17338
rect 321652 17274 321704 17280
rect 321112 16546 321324 16574
rect 320824 4208 320876 4214
rect 320824 4150 320876 4156
rect 320548 3664 320600 3670
rect 320548 3606 320600 3612
rect 321296 3534 321324 16546
rect 322216 15978 322244 84166
rect 322584 57322 322612 84166
rect 322768 69698 322796 84166
rect 322756 69692 322808 69698
rect 322756 69634 322808 69640
rect 322572 57316 322624 57322
rect 322572 57258 322624 57264
rect 323136 55962 323164 84166
rect 323124 55956 323176 55962
rect 323124 55898 323176 55904
rect 322940 54528 322992 54534
rect 322940 54470 322992 54476
rect 322952 16574 322980 54470
rect 323320 31074 323348 84166
rect 323308 31068 323360 31074
rect 323308 31010 323360 31016
rect 322952 16546 323440 16574
rect 322204 15972 322256 15978
rect 322204 15914 322256 15920
rect 322296 4208 322348 4214
rect 322296 4150 322348 4156
rect 321284 3528 321336 3534
rect 320468 3454 321232 3482
rect 321284 3470 321336 3476
rect 321204 480 321232 3454
rect 322308 480 322336 4150
rect 323412 480 323440 16546
rect 323596 4214 323624 93826
rect 323688 54534 323716 96886
rect 323768 96824 323820 96830
rect 323768 96766 323820 96772
rect 323676 54528 323728 54534
rect 323676 54470 323728 54476
rect 323780 4826 323808 96766
rect 323872 29646 323900 96886
rect 324056 96778 324084 97378
rect 323964 96750 324084 96778
rect 323964 82142 323992 96750
rect 324148 93226 324176 100028
rect 324136 93220 324188 93226
rect 324136 93162 324188 93168
rect 323952 82136 324004 82142
rect 323952 82078 324004 82084
rect 324332 53106 324360 100028
rect 324516 84194 324544 100028
rect 324700 97510 324728 100028
rect 324688 97504 324740 97510
rect 324688 97446 324740 97452
rect 324884 84194 324912 100028
rect 325068 96914 325096 100028
rect 324424 84166 324544 84194
rect 324792 84166 324912 84194
rect 324976 96886 325096 96914
rect 324424 72554 324452 84166
rect 324412 72548 324464 72554
rect 324412 72490 324464 72496
rect 324792 68406 324820 84166
rect 324780 68400 324832 68406
rect 324780 68342 324832 68348
rect 324320 53100 324372 53106
rect 324320 53042 324372 53048
rect 324320 32428 324372 32434
rect 324320 32370 324372 32376
rect 323860 29640 323912 29646
rect 323860 29582 323912 29588
rect 324332 16574 324360 32370
rect 324976 28286 325004 96886
rect 325056 96756 325108 96762
rect 325056 96698 325108 96704
rect 324964 28280 325016 28286
rect 324964 28222 325016 28228
rect 324332 16546 324544 16574
rect 323768 4820 323820 4826
rect 323768 4762 323820 4768
rect 323584 4208 323636 4214
rect 323584 4150 323636 4156
rect 324516 480 324544 16546
rect 325068 14550 325096 96698
rect 325252 90438 325280 100028
rect 325240 90432 325292 90438
rect 325240 90374 325292 90380
rect 325436 84194 325464 100028
rect 325620 84194 325648 100028
rect 325804 97782 325832 100028
rect 325792 97776 325844 97782
rect 325792 97718 325844 97724
rect 325988 84194 326016 100028
rect 326172 84194 326200 100028
rect 326356 97866 326384 100028
rect 326356 97838 326476 97866
rect 326344 97708 326396 97714
rect 326344 97650 326396 97656
rect 325344 84166 325464 84194
rect 325528 84166 325648 84194
rect 325896 84166 326016 84194
rect 326080 84166 326200 84194
rect 325344 50454 325372 84166
rect 325332 50448 325384 50454
rect 325332 50390 325384 50396
rect 325528 26926 325556 84166
rect 325896 66910 325924 84166
rect 325884 66904 325936 66910
rect 325884 66846 325936 66852
rect 326080 50386 326108 84166
rect 326356 76634 326384 97650
rect 326448 97306 326476 97838
rect 326436 97300 326488 97306
rect 326436 97242 326488 97248
rect 326540 84194 326568 100028
rect 326724 84194 326752 100028
rect 326908 97442 326936 100028
rect 326896 97436 326948 97442
rect 326896 97378 326948 97384
rect 326448 84166 326568 84194
rect 326632 84166 326752 84194
rect 326344 76628 326396 76634
rect 326344 76570 326396 76576
rect 326068 50380 326120 50386
rect 326068 50322 326120 50328
rect 326448 47666 326476 84166
rect 326436 47660 326488 47666
rect 326436 47602 326488 47608
rect 325516 26920 325568 26926
rect 325516 26862 325568 26868
rect 326632 25566 326660 84166
rect 327092 46306 327120 100028
rect 327276 84194 327304 100028
rect 327460 95946 327488 100028
rect 327448 95940 327500 95946
rect 327448 95882 327500 95888
rect 327644 84194 327672 100028
rect 327828 84194 327856 100028
rect 328012 86290 328040 100028
rect 328000 86284 328052 86290
rect 328000 86226 328052 86232
rect 328196 84194 328224 100028
rect 328380 84194 328408 100028
rect 328564 84862 328592 100028
rect 328552 84856 328604 84862
rect 328552 84798 328604 84804
rect 328748 84194 328776 100028
rect 328932 84194 328960 100028
rect 329116 84194 329144 100028
rect 329300 84194 329328 100028
rect 329484 84194 329512 100028
rect 329668 84194 329696 100028
rect 329852 89010 329880 100028
rect 329840 89004 329892 89010
rect 329840 88946 329892 88952
rect 330036 84194 330064 100028
rect 330220 97238 330248 100028
rect 330208 97232 330260 97238
rect 330208 97174 330260 97180
rect 330404 84194 330432 100028
rect 330588 84194 330616 100028
rect 330772 97714 330800 100028
rect 330760 97708 330812 97714
rect 330760 97650 330812 97656
rect 330956 84194 330984 100028
rect 331140 84194 331168 100028
rect 331324 94518 331352 100028
rect 331220 94512 331272 94518
rect 331220 94454 331272 94460
rect 331312 94512 331364 94518
rect 331312 94454 331364 94460
rect 327184 84166 327304 84194
rect 327552 84166 327672 84194
rect 327736 84166 327856 84194
rect 328104 84166 328224 84194
rect 328288 84166 328408 84194
rect 328656 84166 328776 84194
rect 328840 84166 328960 84194
rect 329024 84166 329144 84194
rect 329208 84166 329328 84194
rect 329392 84166 329512 84194
rect 329576 84166 329696 84194
rect 329944 84166 330064 84194
rect 330312 84166 330432 84194
rect 330496 84166 330616 84194
rect 330864 84166 330984 84194
rect 331048 84166 331168 84194
rect 327184 58682 327212 84166
rect 327552 65550 327580 84166
rect 327540 65544 327592 65550
rect 327540 65486 327592 65492
rect 327172 58676 327224 58682
rect 327172 58618 327224 58624
rect 327080 46300 327132 46306
rect 327080 46242 327132 46248
rect 327080 44872 327132 44878
rect 327080 44814 327132 44820
rect 326620 25560 326672 25566
rect 326620 25502 326672 25508
rect 327092 16574 327120 44814
rect 327736 24138 327764 84166
rect 328104 44946 328132 84166
rect 328092 44940 328144 44946
rect 328092 44882 328144 44888
rect 327724 24132 327776 24138
rect 327724 24074 327776 24080
rect 328288 21418 328316 84166
rect 328460 82136 328512 82142
rect 328460 82078 328512 82084
rect 328276 21412 328328 21418
rect 328276 21354 328328 21360
rect 328472 16574 328500 82078
rect 328656 43518 328684 84166
rect 328840 47598 328868 84166
rect 329024 83502 329052 84166
rect 329012 83496 329064 83502
rect 329012 83438 329064 83444
rect 328828 47592 328880 47598
rect 328828 47534 328880 47540
rect 328644 43512 328696 43518
rect 328644 43454 328696 43460
rect 329208 42158 329236 84166
rect 329196 42152 329248 42158
rect 329196 42094 329248 42100
rect 327092 16546 327856 16574
rect 328472 16546 328960 16574
rect 325056 14544 325108 14550
rect 325056 14486 325108 14492
rect 326712 11756 326764 11762
rect 326712 11698 326764 11704
rect 325608 4208 325660 4214
rect 325608 4150 325660 4156
rect 325620 480 325648 4150
rect 326724 480 326752 11698
rect 327828 480 327856 16546
rect 328932 480 328960 16546
rect 329392 14482 329420 84166
rect 329576 82210 329604 84166
rect 329564 82204 329616 82210
rect 329564 82146 329616 82152
rect 329944 46238 329972 84166
rect 330312 80714 330340 84166
rect 330300 80708 330352 80714
rect 330300 80650 330352 80656
rect 329840 46232 329892 46238
rect 329840 46174 329892 46180
rect 329932 46232 329984 46238
rect 329932 46174 329984 46180
rect 329380 14476 329432 14482
rect 329380 14418 329432 14424
rect 329852 2446 329880 46174
rect 330496 19990 330524 84166
rect 330864 64190 330892 84166
rect 330852 64184 330904 64190
rect 330852 64126 330904 64132
rect 331048 57254 331076 84166
rect 331036 57248 331088 57254
rect 331036 57190 331088 57196
rect 330484 19984 330536 19990
rect 330484 19926 330536 19932
rect 331232 16574 331260 94454
rect 331508 84194 331536 100028
rect 331692 84194 331720 100028
rect 331876 84194 331904 100028
rect 332060 84194 332088 100028
rect 332244 84194 332272 100028
rect 332428 84194 332456 100028
rect 332612 93854 332640 100028
rect 332612 93826 332732 93854
rect 331416 84166 331536 84194
rect 331600 84166 331720 84194
rect 331784 84166 331904 84194
rect 331968 84166 332088 84194
rect 332152 84166 332272 84194
rect 332336 84166 332456 84194
rect 331416 40730 331444 84166
rect 331404 40724 331456 40730
rect 331404 40666 331456 40672
rect 331600 18630 331628 84166
rect 331784 79354 331812 84166
rect 331772 79348 331824 79354
rect 331772 79290 331824 79296
rect 331968 39370 331996 84166
rect 331956 39364 332008 39370
rect 331956 39306 332008 39312
rect 331588 18624 331640 18630
rect 331588 18566 331640 18572
rect 331232 16546 332088 16574
rect 330024 13116 330076 13122
rect 330024 13058 330076 13064
rect 329840 2440 329892 2446
rect 329840 2382 329892 2388
rect 330036 480 330064 13058
rect 332060 3482 332088 16546
rect 332152 6186 332180 84166
rect 332336 77994 332364 84166
rect 332324 77988 332376 77994
rect 332324 77930 332376 77936
rect 332600 72480 332652 72486
rect 332600 72422 332652 72428
rect 332612 16574 332640 72422
rect 332704 62830 332732 93826
rect 332796 68338 332824 100028
rect 332980 97918 333008 100028
rect 332968 97912 333020 97918
rect 332968 97854 333020 97860
rect 333164 84194 333192 100028
rect 333348 84194 333376 100028
rect 333532 91798 333560 100028
rect 333520 91792 333572 91798
rect 333520 91734 333572 91740
rect 333716 84194 333744 100028
rect 333900 84194 333928 100028
rect 334084 93158 334112 100028
rect 334072 93152 334124 93158
rect 334072 93094 334124 93100
rect 334268 84194 334296 100028
rect 334452 84194 334480 100028
rect 334636 97850 334664 100028
rect 334624 97844 334676 97850
rect 334624 97786 334676 97792
rect 334820 84194 334848 100028
rect 335004 84194 335032 100028
rect 335188 84194 335216 100028
rect 335372 96898 335400 100028
rect 335360 96892 335412 96898
rect 335360 96834 335412 96840
rect 335556 84194 335584 100028
rect 335740 96966 335768 100028
rect 335728 96960 335780 96966
rect 335728 96902 335780 96908
rect 335924 84194 335952 100028
rect 336108 84194 336136 100028
rect 336292 90370 336320 100028
rect 336280 90364 336332 90370
rect 336280 90306 336332 90312
rect 336476 84194 336504 100028
rect 336660 84194 336688 100028
rect 336844 84194 336872 100028
rect 337028 84194 337056 100028
rect 337212 84194 337240 100028
rect 338764 97912 338816 97918
rect 338764 97854 338816 97860
rect 337476 97844 337528 97850
rect 337476 97786 337528 97792
rect 337384 96960 337436 96966
rect 337384 96902 337436 96908
rect 333072 84166 333192 84194
rect 333256 84166 333376 84194
rect 333624 84166 333744 84194
rect 333808 84166 333928 84194
rect 334176 84166 334296 84194
rect 334360 84166 334480 84194
rect 334728 84166 334848 84194
rect 334912 84166 335032 84194
rect 335096 84166 335216 84194
rect 335464 84166 335584 84194
rect 335832 84166 335952 84194
rect 336016 84166 336136 84194
rect 336384 84166 336504 84194
rect 336568 84166 336688 84194
rect 336752 84166 336872 84194
rect 336936 84166 337056 84194
rect 337120 84166 337240 84194
rect 333072 82142 333100 84166
rect 333060 82136 333112 82142
rect 333060 82078 333112 82084
rect 332784 68332 332836 68338
rect 332784 68274 332836 68280
rect 332692 62824 332744 62830
rect 332692 62766 332744 62772
rect 333256 17270 333284 84166
rect 333624 37942 333652 84166
rect 333808 44878 333836 84166
rect 333796 44872 333848 44878
rect 333796 44814 333848 44820
rect 333612 37936 333664 37942
rect 333612 37878 333664 37884
rect 334176 36582 334204 84166
rect 334360 55894 334388 84166
rect 334348 55888 334400 55894
rect 334348 55830 334400 55836
rect 334164 36576 334216 36582
rect 334164 36518 334216 36524
rect 333980 35284 334032 35290
rect 333980 35226 334032 35232
rect 333244 17264 333296 17270
rect 333244 17206 333296 17212
rect 333992 16574 334020 35226
rect 334728 33794 334756 84166
rect 334716 33788 334768 33794
rect 334716 33730 334768 33736
rect 332612 16546 333376 16574
rect 333992 16546 334480 16574
rect 332140 6180 332192 6186
rect 332140 6122 332192 6128
rect 332060 3454 332272 3482
rect 331128 2440 331180 2446
rect 331128 2382 331180 2388
rect 331140 480 331168 2382
rect 332244 480 332272 3454
rect 333348 480 333376 16546
rect 334452 480 334480 16546
rect 334912 15910 334940 84166
rect 335096 73846 335124 84166
rect 335084 73840 335136 73846
rect 335084 73782 335136 73788
rect 335360 61532 335412 61538
rect 335360 61474 335412 61480
rect 334900 15904 334952 15910
rect 334900 15846 334952 15852
rect 335372 2650 335400 61474
rect 335464 43450 335492 84166
rect 335832 60042 335860 84166
rect 335820 60036 335872 60042
rect 335820 59978 335872 59984
rect 335452 43444 335504 43450
rect 335452 43386 335504 43392
rect 336016 42090 336044 84166
rect 336004 42084 336056 42090
rect 336004 42026 336056 42032
rect 336384 32434 336412 84166
rect 336372 32428 336424 32434
rect 336372 32370 336424 32376
rect 336568 4826 336596 84166
rect 335544 4820 335596 4826
rect 335544 4762 335596 4768
rect 336556 4820 336608 4826
rect 336556 4762 336608 4768
rect 335360 2644 335412 2650
rect 335360 2586 335412 2592
rect 335556 480 335584 4762
rect 336752 3194 336780 84166
rect 336832 22840 336884 22846
rect 336832 22782 336884 22788
rect 336844 3482 336872 22782
rect 336936 3602 336964 84166
rect 337120 3641 337148 84166
rect 337396 72486 337424 96902
rect 337488 76566 337516 97786
rect 338120 96280 338172 96286
rect 338120 96222 338172 96228
rect 337476 76560 337528 76566
rect 337476 76502 337528 76508
rect 337384 72480 337436 72486
rect 337384 72422 337436 72428
rect 338132 6914 338160 96222
rect 338776 11762 338804 97854
rect 339040 97776 339092 97782
rect 339040 97718 339092 97724
rect 338856 97640 338908 97646
rect 338856 97582 338908 97588
rect 338868 51746 338896 97582
rect 338948 97232 339000 97238
rect 338948 97174 339000 97180
rect 338960 80782 338988 97174
rect 339052 89078 339080 97718
rect 347044 97708 347096 97714
rect 347044 97650 347096 97656
rect 341524 97572 341576 97578
rect 341524 97514 341576 97520
rect 340144 96892 340196 96898
rect 340144 96834 340196 96840
rect 339500 90636 339552 90642
rect 339500 90578 339552 90584
rect 339040 89072 339092 89078
rect 339040 89014 339092 89020
rect 338948 80776 339000 80782
rect 338948 80718 339000 80724
rect 338856 51740 338908 51746
rect 338856 51682 338908 51688
rect 339512 16574 339540 90578
rect 339512 16546 340000 16574
rect 338764 11756 338816 11762
rect 338764 11698 338816 11704
rect 338132 6886 338896 6914
rect 337106 3632 337162 3641
rect 336924 3596 336976 3602
rect 337106 3567 337162 3576
rect 336924 3538 336976 3544
rect 336844 3454 337792 3482
rect 336740 3188 336792 3194
rect 336740 3130 336792 3136
rect 336648 2644 336700 2650
rect 336648 2586 336700 2592
rect 336660 480 336688 2586
rect 337764 480 337792 3454
rect 338868 480 338896 6886
rect 339972 480 340000 16546
rect 340156 13122 340184 96834
rect 340880 91928 340932 91934
rect 340880 91870 340932 91876
rect 340144 13116 340196 13122
rect 340144 13058 340196 13064
rect 340892 3466 340920 91870
rect 340972 80912 341024 80918
rect 340972 80854 341024 80860
rect 340984 16574 341012 80854
rect 340984 16546 341104 16574
rect 340880 3460 340932 3466
rect 340880 3402 340932 3408
rect 341076 480 341104 16546
rect 341536 4894 341564 97514
rect 342904 97504 342956 97510
rect 342904 97446 342956 97452
rect 342260 76764 342312 76770
rect 342260 76706 342312 76712
rect 342272 16574 342300 76706
rect 342272 16546 342852 16574
rect 341524 4888 341576 4894
rect 341524 4830 341576 4836
rect 342824 3482 342852 16546
rect 342916 6254 342944 97446
rect 345664 97436 345716 97442
rect 345664 97378 345716 97384
rect 345020 93356 345072 93362
rect 345020 93298 345072 93304
rect 345032 16574 345060 93298
rect 345032 16546 345520 16574
rect 344376 10328 344428 10334
rect 344376 10270 344428 10276
rect 342904 6248 342956 6254
rect 342904 6190 342956 6196
rect 342168 3460 342220 3466
rect 342168 3402 342220 3408
rect 342260 3460 342312 3466
rect 342824 3454 343312 3482
rect 342260 3402 342312 3408
rect 342180 480 342208 3402
rect 342272 3194 342300 3402
rect 342260 3188 342312 3194
rect 342260 3130 342312 3136
rect 343284 480 343312 3454
rect 344388 480 344416 10270
rect 345492 480 345520 16546
rect 345676 7614 345704 97378
rect 346400 93424 346452 93430
rect 346400 93366 346452 93372
rect 345664 7608 345716 7614
rect 345664 7550 345716 7556
rect 346412 3482 346440 93366
rect 346492 40860 346544 40866
rect 346492 40802 346544 40808
rect 346504 4214 346532 40802
rect 347056 10334 347084 97650
rect 349804 97368 349856 97374
rect 349804 97310 349856 97316
rect 349816 91934 349844 97310
rect 349804 91928 349856 91934
rect 349804 91870 349856 91876
rect 347780 89276 347832 89282
rect 347780 89218 347832 89224
rect 347792 16574 347820 89218
rect 351920 87848 351972 87854
rect 351920 87790 351972 87796
rect 350540 82340 350592 82346
rect 350540 82282 350592 82288
rect 349160 75336 349212 75342
rect 349160 75278 349212 75284
rect 349172 16574 349200 75278
rect 350552 16574 350580 82282
rect 347792 16546 348832 16574
rect 349172 16546 349936 16574
rect 350552 16546 351040 16574
rect 347044 10328 347096 10334
rect 347044 10270 347096 10276
rect 346492 4208 346544 4214
rect 346492 4150 346544 4156
rect 347688 4208 347740 4214
rect 347688 4150 347740 4156
rect 346412 3454 346624 3482
rect 346596 480 346624 3454
rect 347700 480 347728 4150
rect 348804 480 348832 16546
rect 349908 480 349936 16546
rect 351012 480 351040 16546
rect 351932 3482 351960 87790
rect 352012 79552 352064 79558
rect 352012 79494 352064 79500
rect 352024 4214 352052 79494
rect 353300 33924 353352 33930
rect 353300 33866 353352 33872
rect 353312 6914 353340 33866
rect 353956 9654 353984 102031
rect 354048 23458 354076 105567
rect 354140 35902 354168 109103
rect 354232 49706 354260 112639
rect 354324 62082 354352 116175
rect 354416 75886 354444 119711
rect 354508 88330 354536 123247
rect 354600 102134 354628 126783
rect 580172 114504 580224 114510
rect 580170 114472 580172 114481
rect 580224 114472 580226 114481
rect 580170 114407 580226 114416
rect 354588 102128 354640 102134
rect 354588 102070 354640 102076
rect 579988 102128 580040 102134
rect 579988 102070 580040 102076
rect 580000 101289 580028 102070
rect 579986 101280 580042 101289
rect 579986 101215 580042 101224
rect 475384 97300 475436 97306
rect 475384 97242 475436 97248
rect 354680 96212 354732 96218
rect 354680 96154 354732 96160
rect 354496 88324 354548 88330
rect 354496 88266 354548 88272
rect 354404 75880 354456 75886
rect 354404 75822 354456 75828
rect 354312 62076 354364 62082
rect 354312 62018 354364 62024
rect 354220 49700 354272 49706
rect 354220 49642 354272 49648
rect 354128 35896 354180 35902
rect 354128 35838 354180 35844
rect 354036 23452 354088 23458
rect 354036 23394 354088 23400
rect 354692 16574 354720 96154
rect 390560 96144 390612 96150
rect 390560 96086 390612 96092
rect 357440 94784 357492 94790
rect 357440 94726 357492 94732
rect 356060 72684 356112 72690
rect 356060 72626 356112 72632
rect 356072 16574 356100 72626
rect 354692 16546 355456 16574
rect 356072 16546 356560 16574
rect 353944 9648 353996 9654
rect 353944 9590 353996 9596
rect 353312 6886 354352 6914
rect 352012 4208 352064 4214
rect 352012 4150 352064 4156
rect 353208 4208 353260 4214
rect 353208 4150 353260 4156
rect 351932 3454 352144 3482
rect 352116 480 352144 3454
rect 353220 480 353248 4150
rect 354324 480 354352 6886
rect 355428 480 355456 16546
rect 356532 480 356560 16546
rect 357452 3194 357480 94726
rect 387800 93288 387852 93294
rect 387800 93230 387852 93236
rect 361580 92064 361632 92070
rect 361580 92006 361632 92012
rect 358820 78192 358872 78198
rect 358820 78134 358872 78140
rect 358832 16574 358860 78134
rect 360200 39500 360252 39506
rect 360200 39442 360252 39448
rect 360212 16574 360240 39442
rect 361592 16574 361620 92006
rect 386420 91996 386472 92002
rect 386420 91938 386472 91944
rect 362960 90568 363012 90574
rect 362960 90510 363012 90516
rect 358832 16546 359872 16574
rect 360212 16546 360976 16574
rect 361592 16546 362080 16574
rect 357624 8968 357676 8974
rect 357624 8910 357676 8916
rect 357440 3188 357492 3194
rect 357440 3130 357492 3136
rect 357636 480 357664 8910
rect 358728 3188 358780 3194
rect 358728 3130 358780 3136
rect 358740 480 358768 3130
rect 359844 480 359872 16546
rect 360948 480 360976 16546
rect 362052 480 362080 16546
rect 362972 3482 363000 90510
rect 364340 90500 364392 90506
rect 364340 90442 364392 90448
rect 363052 67040 363104 67046
rect 363052 66982 363104 66988
rect 363064 4214 363092 66982
rect 364352 16574 364380 90442
rect 371240 89208 371292 89214
rect 371240 89150 371292 89156
rect 368480 86488 368532 86494
rect 368480 86430 368532 86436
rect 365720 61464 365772 61470
rect 365720 61406 365772 61412
rect 365732 16574 365760 61406
rect 367100 38004 367152 38010
rect 367100 37946 367152 37952
rect 367112 16574 367140 37946
rect 364352 16546 365392 16574
rect 365732 16546 366496 16574
rect 367112 16546 367600 16574
rect 363052 4208 363104 4214
rect 363052 4150 363104 4156
rect 364248 4208 364300 4214
rect 364248 4150 364300 4156
rect 362972 3454 363184 3482
rect 363156 480 363184 3454
rect 364260 480 364288 4150
rect 365364 480 365392 16546
rect 366468 480 366496 16546
rect 367572 480 367600 16546
rect 368492 3482 368520 86430
rect 368572 73976 368624 73982
rect 368572 73918 368624 73924
rect 368584 4214 368612 73918
rect 369860 36644 369912 36650
rect 369860 36586 369912 36592
rect 369872 16574 369900 36586
rect 371252 16574 371280 89150
rect 374000 87780 374052 87786
rect 374000 87722 374052 87728
rect 372620 76696 372672 76702
rect 372620 76638 372672 76644
rect 372632 16574 372660 76638
rect 369872 16546 370912 16574
rect 371252 16546 372016 16574
rect 372632 16546 373120 16574
rect 368572 4208 368624 4214
rect 368572 4150 368624 4156
rect 369768 4208 369820 4214
rect 369768 4150 369820 4156
rect 368492 3454 368704 3482
rect 368676 480 368704 3454
rect 369780 480 369808 4150
rect 370884 480 370912 16546
rect 371988 480 372016 16546
rect 373092 480 373120 16546
rect 374012 3194 374040 87722
rect 385040 86420 385092 86426
rect 385040 86362 385092 86368
rect 378140 85060 378192 85066
rect 378140 85002 378192 85008
rect 375380 49088 375432 49094
rect 375380 49030 375432 49036
rect 375392 16574 375420 49030
rect 376760 35216 376812 35222
rect 376760 35158 376812 35164
rect 376772 16574 376800 35158
rect 378152 16574 378180 85002
rect 380900 83700 380952 83706
rect 380900 83642 380952 83648
rect 379520 58812 379572 58818
rect 379520 58754 379572 58760
rect 375392 16546 376432 16574
rect 376772 16546 377536 16574
rect 378152 16546 378640 16574
rect 374184 7676 374236 7682
rect 374184 7618 374236 7624
rect 374000 3188 374052 3194
rect 374000 3130 374052 3136
rect 374196 480 374224 7618
rect 375288 3188 375340 3194
rect 375288 3130 375340 3136
rect 375300 480 375328 3130
rect 376404 480 376432 16546
rect 377508 480 377536 16546
rect 378612 480 378640 16546
rect 379532 3482 379560 58754
rect 380912 16574 380940 83642
rect 382280 57384 382332 57390
rect 382280 57326 382332 57332
rect 382292 16574 382320 57326
rect 383660 22772 383712 22778
rect 383660 22714 383712 22720
rect 383672 16574 383700 22714
rect 380912 16546 381952 16574
rect 382292 16546 383056 16574
rect 383672 16546 384160 16574
rect 379612 11824 379664 11830
rect 379612 11766 379664 11772
rect 379624 4214 379652 11766
rect 379612 4208 379664 4214
rect 379612 4150 379664 4156
rect 380808 4208 380860 4214
rect 380808 4150 380860 4156
rect 379532 3454 379744 3482
rect 379716 480 379744 3454
rect 380820 480 380848 4150
rect 381924 480 381952 16546
rect 383028 480 383056 16546
rect 384132 480 384160 16546
rect 385052 3194 385080 86362
rect 385132 80844 385184 80850
rect 385132 80786 385184 80792
rect 385144 16574 385172 80786
rect 386432 16574 386460 91938
rect 387812 16574 387840 93230
rect 389180 87712 389232 87718
rect 389180 87654 389232 87660
rect 389192 16574 389220 87654
rect 385144 16546 385264 16574
rect 386432 16546 387472 16574
rect 387812 16546 388576 16574
rect 389192 16546 389680 16574
rect 385040 3188 385092 3194
rect 385040 3130 385092 3136
rect 385236 480 385264 16546
rect 386328 3188 386380 3194
rect 386328 3130 386380 3136
rect 386340 480 386368 3130
rect 387444 480 387472 16546
rect 388548 480 388576 16546
rect 389652 480 389680 16546
rect 390572 3194 390600 96086
rect 434720 96076 434772 96082
rect 434720 96018 434772 96024
rect 402980 94716 403032 94722
rect 402980 94658 403032 94664
rect 394700 82272 394752 82278
rect 394700 82214 394752 82220
rect 391940 72616 391992 72622
rect 391940 72558 391992 72564
rect 390652 32496 390704 32502
rect 390652 32438 390704 32444
rect 390664 16574 390692 32438
rect 391952 16574 391980 72558
rect 394712 16574 394740 82214
rect 397460 71188 397512 71194
rect 397460 71130 397512 71136
rect 396080 65680 396132 65686
rect 396080 65622 396132 65628
rect 390664 16546 390784 16574
rect 391952 16546 392992 16574
rect 394712 16546 395200 16574
rect 390560 3188 390612 3194
rect 390560 3130 390612 3136
rect 390756 480 390784 16546
rect 391848 3188 391900 3194
rect 391848 3130 391900 3136
rect 391860 480 391888 3130
rect 392964 480 392992 16546
rect 394056 13184 394108 13190
rect 394056 13126 394108 13132
rect 394068 480 394096 13126
rect 395172 480 395200 16546
rect 396092 3194 396120 65622
rect 396172 56024 396224 56030
rect 396172 55966 396224 55972
rect 396184 16574 396212 55966
rect 397472 16574 397500 71130
rect 401600 69828 401652 69834
rect 401600 69770 401652 69776
rect 398840 51808 398892 51814
rect 398840 51750 398892 51756
rect 398852 16574 398880 51750
rect 396184 16546 396304 16574
rect 397472 16546 398512 16574
rect 398852 16546 399616 16574
rect 396080 3188 396132 3194
rect 396080 3130 396132 3136
rect 396276 480 396304 16546
rect 397368 3188 397420 3194
rect 397368 3130 397420 3136
rect 397380 480 397408 3130
rect 398484 480 398512 16546
rect 399588 480 399616 16546
rect 400680 10396 400732 10402
rect 400680 10338 400732 10344
rect 400692 480 400720 10338
rect 401612 3482 401640 69770
rect 401692 53168 401744 53174
rect 401692 53110 401744 53116
rect 401704 4214 401732 53110
rect 402992 16574 403020 94658
rect 420920 94648 420972 94654
rect 420920 94590 420972 94596
rect 411260 89140 411312 89146
rect 411260 89082 411312 89088
rect 404360 86352 404412 86358
rect 404360 86294 404412 86300
rect 404372 16574 404400 86294
rect 407120 79484 407172 79490
rect 407120 79426 407172 79432
rect 405740 75268 405792 75274
rect 405740 75210 405792 75216
rect 405752 16574 405780 75210
rect 402992 16546 404032 16574
rect 404372 16546 405136 16574
rect 405752 16546 406240 16574
rect 401692 4208 401744 4214
rect 401692 4150 401744 4156
rect 402888 4208 402940 4214
rect 402888 4150 402940 4156
rect 401612 3454 401824 3482
rect 401796 480 401824 3454
rect 402900 480 402928 4150
rect 404004 480 404032 16546
rect 405108 480 405136 16546
rect 406212 480 406240 16546
rect 407132 3194 407160 79426
rect 409880 49020 409932 49026
rect 409880 48962 409932 48968
rect 407212 40792 407264 40798
rect 407212 40734 407264 40740
rect 407224 16574 407252 40734
rect 408500 31136 408552 31142
rect 408500 31078 408552 31084
rect 408512 16574 408540 31078
rect 409892 16574 409920 48962
rect 411272 16574 411300 89082
rect 414020 87644 414072 87650
rect 414020 87586 414072 87592
rect 412640 84992 412692 84998
rect 412640 84934 412692 84940
rect 407224 16546 407344 16574
rect 408512 16546 409552 16574
rect 409892 16546 410656 16574
rect 411272 16546 411760 16574
rect 407120 3188 407172 3194
rect 407120 3130 407172 3136
rect 407316 480 407344 16546
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 408420 480 408448 3130
rect 409524 480 409552 16546
rect 410628 480 410656 16546
rect 411732 480 411760 16546
rect 412652 3482 412680 84934
rect 412732 62960 412784 62966
rect 412732 62902 412784 62908
rect 412744 4214 412772 62902
rect 414032 16574 414060 87586
rect 418160 79416 418212 79422
rect 418160 79358 418212 79364
rect 416780 39432 416832 39438
rect 416780 39374 416832 39380
rect 415400 29708 415452 29714
rect 415400 29650 415452 29656
rect 415412 16574 415440 29650
rect 416792 16574 416820 39374
rect 414032 16546 415072 16574
rect 415412 16546 416176 16574
rect 416792 16546 417280 16574
rect 412732 4208 412784 4214
rect 412732 4150 412784 4156
rect 413928 4208 413980 4214
rect 413928 4150 413980 4156
rect 412652 3454 412864 3482
rect 412836 480 412864 3454
rect 413940 480 413968 4150
rect 415044 480 415072 16546
rect 416148 480 416176 16546
rect 417252 480 417280 16546
rect 418172 3262 418200 79358
rect 418252 78124 418304 78130
rect 418252 78066 418304 78072
rect 418264 16574 418292 78066
rect 419540 60172 419592 60178
rect 419540 60114 419592 60120
rect 419552 16574 419580 60114
rect 420932 16574 420960 94590
rect 427820 84924 427872 84930
rect 427820 84866 427872 84872
rect 423680 75200 423732 75206
rect 423680 75142 423732 75148
rect 422300 54596 422352 54602
rect 422300 54538 422352 54544
rect 422312 16574 422340 54538
rect 418264 16546 418384 16574
rect 419552 16546 420592 16574
rect 420932 16546 421696 16574
rect 422312 16546 422800 16574
rect 418160 3256 418212 3262
rect 418160 3198 418212 3204
rect 418356 480 418384 16546
rect 419448 3256 419500 3262
rect 419448 3198 419500 3204
rect 419460 480 419488 3198
rect 420564 480 420592 16546
rect 421668 480 421696 16546
rect 422772 480 422800 16546
rect 423692 3262 423720 75142
rect 426440 64320 426492 64326
rect 426440 64262 426492 64268
rect 423772 33856 423824 33862
rect 423772 33798 423824 33804
rect 423784 16574 423812 33798
rect 425060 28348 425112 28354
rect 425060 28290 425112 28296
rect 425072 16574 425100 28290
rect 426452 16574 426480 64262
rect 427832 16574 427860 84866
rect 430580 68468 430632 68474
rect 430580 68410 430632 68416
rect 429292 26988 429344 26994
rect 429292 26930 429344 26936
rect 429304 16574 429332 26930
rect 430592 16574 430620 68410
rect 431960 25628 432012 25634
rect 431960 25570 432012 25576
rect 431972 16574 432000 25570
rect 423784 16546 423904 16574
rect 425072 16546 426112 16574
rect 426452 16546 427216 16574
rect 427832 16546 428320 16574
rect 429304 16546 429424 16574
rect 430592 16546 431632 16574
rect 431972 16546 432736 16574
rect 423680 3256 423732 3262
rect 423680 3198 423732 3204
rect 423876 480 423904 16546
rect 424968 3256 425020 3262
rect 424968 3198 425020 3204
rect 424980 480 425008 3198
rect 426084 480 426112 16546
rect 427188 480 427216 16546
rect 428292 480 428320 16546
rect 429396 480 429424 16546
rect 430488 3188 430540 3194
rect 430488 3130 430540 3136
rect 430500 480 430528 3130
rect 431604 480 431632 16546
rect 432708 480 432736 16546
rect 434732 3398 434760 96018
rect 467840 91928 467892 91934
rect 467840 91870 467892 91876
rect 454040 91860 454092 91866
rect 454040 91802 454092 91808
rect 440332 83632 440384 83638
rect 440332 83574 440384 83580
rect 437480 76628 437532 76634
rect 437480 76570 437532 76576
rect 434812 66972 434864 66978
rect 434812 66914 434864 66920
rect 434824 16574 434852 66914
rect 437492 16574 437520 76570
rect 438860 71120 438912 71126
rect 438860 71062 438912 71068
rect 438872 16574 438900 71062
rect 434824 16546 434944 16574
rect 437492 16546 438256 16574
rect 438872 16546 439360 16574
rect 434720 3392 434772 3398
rect 434720 3334 434772 3340
rect 433800 3324 433852 3330
rect 433800 3266 433852 3272
rect 433812 480 433840 3266
rect 434916 480 434944 16546
rect 436008 3392 436060 3398
rect 436008 3334 436060 3340
rect 436020 480 436048 3334
rect 437112 3324 437164 3330
rect 437112 3266 437164 3272
rect 437124 480 437152 3266
rect 438228 480 438256 16546
rect 439332 480 439360 16546
rect 440344 3398 440372 83574
rect 441620 78056 441672 78062
rect 441620 77998 441672 78004
rect 441632 16574 441660 77998
rect 444380 65612 444432 65618
rect 444380 65554 444432 65560
rect 444392 16574 444420 65554
rect 447140 64252 447192 64258
rect 447140 64194 447192 64200
rect 445852 24200 445904 24206
rect 445852 24142 445904 24148
rect 445864 16574 445892 24142
rect 447152 16574 447180 64194
rect 451280 62892 451332 62898
rect 451280 62834 451332 62840
rect 448520 21480 448572 21486
rect 448520 21422 448572 21428
rect 448532 16574 448560 21422
rect 441632 16546 442672 16574
rect 444392 16546 444880 16574
rect 445864 16546 445984 16574
rect 447152 16546 448192 16574
rect 448532 16546 449296 16574
rect 440424 4140 440476 4146
rect 440424 4082 440476 4088
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 440436 480 440464 4082
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 443736 4072 443788 4078
rect 443736 4014 443788 4020
rect 443748 480 443776 4014
rect 444852 480 444880 16546
rect 445956 480 445984 16546
rect 447048 4004 447100 4010
rect 447048 3946 447100 3952
rect 447060 480 447088 3946
rect 448164 480 448192 16546
rect 449268 480 449296 16546
rect 450360 3936 450412 3942
rect 450360 3878 450412 3884
rect 450372 480 450400 3878
rect 451292 3482 451320 62834
rect 454052 16574 454080 91802
rect 462412 83564 462464 83570
rect 462412 83506 462464 83512
rect 456892 71052 456944 71058
rect 456892 70994 456944 71000
rect 455420 61396 455472 61402
rect 455420 61338 455472 61344
rect 455432 16574 455460 61338
rect 454052 16546 454816 16574
rect 455432 16546 455920 16574
rect 451372 14544 451424 14550
rect 451372 14486 451424 14492
rect 451384 4078 451412 14486
rect 451372 4072 451424 4078
rect 451372 4014 451424 4020
rect 452568 4072 452620 4078
rect 452568 4014 452620 4020
rect 451292 3454 451504 3482
rect 451476 480 451504 3454
rect 452580 480 452608 4014
rect 453672 4004 453724 4010
rect 453672 3946 453724 3952
rect 453684 480 453712 3946
rect 454788 480 454816 16546
rect 455892 480 455920 16546
rect 456904 3398 456932 70994
rect 460940 69760 460992 69766
rect 460940 69702 460992 69708
rect 458180 20052 458232 20058
rect 458180 19994 458232 20000
rect 458192 16574 458220 19994
rect 460952 16574 460980 69702
rect 462424 16574 462452 83506
rect 463700 60104 463752 60110
rect 463700 60046 463752 60052
rect 463712 16574 463740 60046
rect 465080 18692 465132 18698
rect 465080 18634 465132 18640
rect 465092 16574 465120 18634
rect 458192 16546 459232 16574
rect 460952 16546 461440 16574
rect 462424 16546 462544 16574
rect 463712 16546 464752 16574
rect 465092 16546 465856 16574
rect 456984 3800 457036 3806
rect 456984 3742 457036 3748
rect 456892 3392 456944 3398
rect 456892 3334 456944 3340
rect 456996 480 457024 3742
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 460296 3732 460348 3738
rect 460296 3674 460348 3680
rect 460308 480 460336 3674
rect 461412 480 461440 16546
rect 462516 480 462544 16546
rect 463608 3664 463660 3670
rect 463608 3606 463660 3612
rect 463620 480 463648 3606
rect 464724 480 464752 16546
rect 465828 480 465856 16546
rect 466920 3528 466972 3534
rect 466920 3470 466972 3476
rect 467852 3482 467880 91870
rect 467932 73908 467984 73914
rect 467932 73850 467984 73856
rect 467944 3670 467972 73850
rect 471980 58744 472032 58750
rect 471980 58686 472032 58692
rect 470600 51740 470652 51746
rect 470600 51682 470652 51688
rect 469220 17332 469272 17338
rect 469220 17274 469272 17280
rect 469232 16574 469260 17274
rect 470612 16574 470640 51682
rect 471992 16574 472020 58686
rect 474740 57316 474792 57322
rect 474740 57258 474792 57264
rect 474752 16574 474780 57258
rect 469232 16546 470272 16574
rect 470612 16546 471376 16574
rect 471992 16546 472480 16574
rect 474752 16546 475332 16574
rect 467932 3664 467984 3670
rect 467932 3606 467984 3612
rect 469128 3664 469180 3670
rect 469128 3606 469180 3612
rect 466932 480 466960 3470
rect 467852 3454 468064 3482
rect 468036 480 468064 3454
rect 469140 480 469168 3606
rect 470244 480 470272 16546
rect 471348 480 471376 16546
rect 472452 480 472480 16546
rect 473544 15972 473596 15978
rect 473544 15914 473596 15920
rect 473556 480 473584 15914
rect 474648 4888 474700 4894
rect 474648 4830 474700 4836
rect 474660 480 474688 4830
rect 475304 3482 475332 16546
rect 475396 4894 475424 97242
rect 477500 96008 477552 96014
rect 477500 95950 477552 95956
rect 476120 69692 476172 69698
rect 476120 69634 476172 69640
rect 476132 16574 476160 69634
rect 477512 16574 477540 95950
rect 503720 95940 503772 95946
rect 503720 95882 503772 95888
rect 480260 94580 480312 94586
rect 480260 94522 480312 94528
rect 478880 55956 478932 55962
rect 478880 55898 478932 55904
rect 476132 16546 476896 16574
rect 477512 16546 478000 16574
rect 475384 4888 475436 4894
rect 475384 4830 475436 4836
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 476868 480 476896 16546
rect 477972 480 478000 16546
rect 478892 3482 478920 55898
rect 478972 31068 479024 31074
rect 478972 31010 479024 31016
rect 478984 3670 479012 31010
rect 480272 16574 480300 94522
rect 484400 93220 484452 93226
rect 484400 93162 484452 93168
rect 481640 54528 481692 54534
rect 481640 54470 481692 54476
rect 481652 16574 481680 54470
rect 483020 29640 483072 29646
rect 483020 29582 483072 29588
rect 483032 16574 483060 29582
rect 480272 16546 481312 16574
rect 481652 16546 482416 16574
rect 483032 16546 483520 16574
rect 478972 3664 479024 3670
rect 478972 3606 479024 3612
rect 480168 3664 480220 3670
rect 480168 3606 480220 3612
rect 478892 3454 479104 3482
rect 479076 480 479104 3454
rect 480180 480 480208 3606
rect 481284 480 481312 16546
rect 482388 480 482416 16546
rect 483492 480 483520 16546
rect 484412 3482 484440 93162
rect 489920 90432 489972 90438
rect 489920 90374 489972 90380
rect 485780 72548 485832 72554
rect 485780 72490 485832 72496
rect 484492 53100 484544 53106
rect 484492 53042 484544 53048
rect 484504 3670 484532 53042
rect 485792 16574 485820 72490
rect 488540 68400 488592 68406
rect 488540 68342 488592 68348
rect 488552 16574 488580 68342
rect 485792 16546 486832 16574
rect 488552 16546 489040 16574
rect 484492 3664 484544 3670
rect 484492 3606 484544 3612
rect 485688 3664 485740 3670
rect 485688 3606 485740 3612
rect 484412 3454 484624 3482
rect 484596 480 484624 3454
rect 485700 480 485728 3606
rect 486804 480 486832 16546
rect 487896 6248 487948 6254
rect 487896 6190 487948 6196
rect 487908 480 487936 6190
rect 489012 480 489040 16546
rect 489932 3534 489960 90374
rect 494060 89072 494112 89078
rect 494060 89014 494112 89020
rect 491300 50448 491352 50454
rect 491300 50390 491352 50396
rect 490012 28280 490064 28286
rect 490012 28222 490064 28228
rect 490024 16574 490052 28222
rect 491312 16574 491340 50390
rect 492680 26920 492732 26926
rect 492680 26862 492732 26868
rect 492692 16574 492720 26862
rect 494072 16574 494100 89014
rect 495440 66904 495492 66910
rect 495440 66846 495492 66852
rect 490024 16546 490144 16574
rect 491312 16546 492352 16574
rect 492692 16546 493456 16574
rect 494072 16546 494560 16574
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490116 480 490144 16546
rect 491208 3528 491260 3534
rect 491208 3470 491260 3476
rect 491220 480 491248 3470
rect 492324 480 492352 16546
rect 493428 480 493456 16546
rect 494532 480 494560 16546
rect 495452 3482 495480 66846
rect 502340 58676 502392 58682
rect 502340 58618 502392 58624
rect 495532 50380 495584 50386
rect 495532 50322 495584 50328
rect 495544 3670 495572 50322
rect 498200 47660 498252 47666
rect 498200 47602 498252 47608
rect 498212 16574 498240 47602
rect 500960 46300 501012 46306
rect 500960 46242 501012 46248
rect 499580 25560 499632 25566
rect 499580 25502 499632 25508
rect 499592 16574 499620 25502
rect 498212 16546 498976 16574
rect 499592 16546 500080 16574
rect 497832 4888 497884 4894
rect 497832 4830 497884 4836
rect 495532 3664 495584 3670
rect 495532 3606 495584 3612
rect 496728 3664 496780 3670
rect 496728 3606 496780 3612
rect 495452 3454 495664 3482
rect 495636 480 495664 3454
rect 496740 480 496768 3606
rect 497844 480 497872 4830
rect 498948 480 498976 16546
rect 500052 480 500080 16546
rect 500972 3534 501000 46242
rect 502352 16574 502380 58618
rect 503732 16574 503760 95882
rect 527180 94512 527232 94518
rect 527180 94454 527232 94460
rect 517520 89004 517572 89010
rect 517520 88946 517572 88952
rect 506480 86284 506532 86290
rect 506480 86226 506532 86232
rect 505100 65544 505152 65550
rect 505100 65486 505152 65492
rect 505112 16574 505140 65486
rect 502352 16546 503392 16574
rect 503732 16546 504496 16574
rect 505112 16546 505600 16574
rect 501144 7608 501196 7614
rect 501144 7550 501196 7556
rect 500960 3528 501012 3534
rect 500960 3470 501012 3476
rect 501156 480 501184 7550
rect 502248 3528 502300 3534
rect 502248 3470 502300 3476
rect 502260 480 502288 3470
rect 503364 480 503392 16546
rect 504468 480 504496 16546
rect 505572 480 505600 16546
rect 506492 3534 506520 86226
rect 510620 84856 510672 84862
rect 510620 84798 510672 84804
rect 507860 44940 507912 44946
rect 507860 44882 507912 44888
rect 506572 24132 506624 24138
rect 506572 24074 506624 24080
rect 506584 16574 506612 24074
rect 507872 16574 507900 44882
rect 509240 21412 509292 21418
rect 509240 21354 509292 21360
rect 509252 16574 509280 21354
rect 510632 16574 510660 84798
rect 513380 83496 513432 83502
rect 513380 83438 513432 83444
rect 512000 47592 512052 47598
rect 512000 47534 512052 47540
rect 506584 16546 506704 16574
rect 507872 16546 508912 16574
rect 509252 16546 510016 16574
rect 510632 16546 511120 16574
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506676 480 506704 16546
rect 507768 3528 507820 3534
rect 507768 3470 507820 3476
rect 507780 480 507808 3470
rect 508884 480 508912 16546
rect 509988 480 510016 16546
rect 511092 480 511120 16546
rect 512012 3534 512040 47534
rect 512092 43512 512144 43518
rect 512092 43454 512144 43460
rect 512104 16574 512132 43454
rect 513392 16574 513420 83438
rect 514760 42152 514812 42158
rect 514760 42094 514812 42100
rect 514772 16574 514800 42094
rect 512104 16546 512224 16574
rect 513392 16546 514432 16574
rect 514772 16546 515536 16574
rect 512000 3528 512052 3534
rect 512000 3470 512052 3476
rect 512196 480 512224 16546
rect 513288 3528 513340 3534
rect 513288 3470 513340 3476
rect 513300 480 513328 3470
rect 514404 480 514432 16546
rect 515508 480 515536 16546
rect 516600 14476 516652 14482
rect 516600 14418 516652 14424
rect 516612 480 516640 14418
rect 517532 3534 517560 88946
rect 517612 82204 517664 82210
rect 517612 82146 517664 82152
rect 517624 16574 517652 82146
rect 520280 80776 520332 80782
rect 520280 80718 520332 80724
rect 518900 46232 518952 46238
rect 518900 46174 518952 46180
rect 518912 16574 518940 46174
rect 520292 16574 520320 80718
rect 521660 80708 521712 80714
rect 521660 80650 521712 80656
rect 521672 16574 521700 80650
rect 524420 64184 524472 64190
rect 524420 64126 524472 64132
rect 523040 19984 523092 19990
rect 523040 19926 523092 19932
rect 517624 16546 517744 16574
rect 518912 16546 519952 16574
rect 520292 16546 521056 16574
rect 521672 16546 522160 16574
rect 517520 3528 517572 3534
rect 517520 3470 517572 3476
rect 517716 480 517744 16546
rect 518808 3528 518860 3534
rect 518808 3470 518860 3476
rect 518820 480 518848 3470
rect 519924 480 519952 16546
rect 521028 480 521056 16546
rect 522132 480 522160 16546
rect 523052 3482 523080 19926
rect 524432 16574 524460 64126
rect 525800 57248 525852 57254
rect 525800 57190 525852 57196
rect 525812 16574 525840 57190
rect 527192 16574 527220 94454
rect 543740 93152 543792 93158
rect 543740 93094 543792 93100
rect 539600 91792 539652 91798
rect 539600 91734 539652 91740
rect 538220 82136 538272 82142
rect 538220 82078 538272 82084
rect 529940 79348 529992 79354
rect 529940 79290 529992 79296
rect 528560 40724 528612 40730
rect 528560 40666 528612 40672
rect 524432 16546 525472 16574
rect 525812 16546 526576 16574
rect 527192 16546 527680 16574
rect 523132 10328 523184 10334
rect 523132 10270 523184 10276
rect 523144 3670 523172 10270
rect 523132 3664 523184 3670
rect 523132 3606 523184 3612
rect 524328 3664 524380 3670
rect 524328 3606 524380 3612
rect 523052 3454 523264 3482
rect 523236 480 523264 3454
rect 524340 480 524368 3606
rect 525444 480 525472 16546
rect 526548 480 526576 16546
rect 527652 480 527680 16546
rect 528572 3482 528600 40666
rect 528652 18624 528704 18630
rect 528652 18566 528704 18572
rect 528664 3670 528692 18566
rect 529952 16574 529980 79290
rect 534080 77988 534132 77994
rect 534080 77930 534132 77936
rect 531320 39364 531372 39370
rect 531320 39306 531372 39312
rect 531332 16574 531360 39306
rect 529952 16546 530992 16574
rect 531332 16546 532096 16574
rect 528652 3664 528704 3670
rect 528652 3606 528704 3612
rect 529848 3664 529900 3670
rect 529848 3606 529900 3612
rect 528572 3454 528784 3482
rect 528756 480 528784 3454
rect 529860 480 529888 3606
rect 530964 480 530992 16546
rect 532068 480 532096 16546
rect 533160 6180 533212 6186
rect 533160 6122 533212 6128
rect 533172 480 533200 6122
rect 534092 3482 534120 77930
rect 535460 68332 535512 68338
rect 535460 68274 535512 68280
rect 534172 62824 534224 62830
rect 534172 62766 534224 62772
rect 534184 3670 534212 62766
rect 535472 16574 535500 68274
rect 538232 16574 538260 82078
rect 535472 16546 536512 16574
rect 538232 16546 538720 16574
rect 534172 3664 534224 3670
rect 534172 3606 534224 3612
rect 535368 3664 535420 3670
rect 535368 3606 535420 3612
rect 534092 3454 534304 3482
rect 534276 480 534304 3454
rect 535380 480 535408 3606
rect 536484 480 536512 16546
rect 537576 11756 537628 11762
rect 537576 11698 537628 11704
rect 537588 480 537616 11698
rect 538692 480 538720 16546
rect 539612 1290 539640 91734
rect 542360 44872 542412 44878
rect 542360 44814 542412 44820
rect 540980 37936 541032 37942
rect 540980 37878 541032 37884
rect 539692 17264 539744 17270
rect 539692 17206 539744 17212
rect 539704 16574 539732 17206
rect 540992 16574 541020 37878
rect 542372 16574 542400 44814
rect 543752 16574 543780 93094
rect 556160 90364 556212 90370
rect 556160 90306 556212 90312
rect 546500 76560 546552 76566
rect 546500 76502 546552 76508
rect 545120 55888 545172 55894
rect 545120 55830 545172 55836
rect 539704 16546 539824 16574
rect 540992 16546 542032 16574
rect 542372 16546 543136 16574
rect 543752 16546 544240 16574
rect 539600 1284 539652 1290
rect 539600 1226 539652 1232
rect 539796 480 539824 16546
rect 540888 1284 540940 1290
rect 540888 1226 540940 1232
rect 540900 480 540928 1226
rect 542004 480 542032 16546
rect 543108 480 543136 16546
rect 544212 480 544240 16546
rect 545132 1290 545160 55830
rect 545212 36576 545264 36582
rect 545212 36518 545264 36524
rect 545224 16574 545252 36518
rect 546512 16574 546540 76502
rect 549904 73840 549956 73846
rect 549904 73782 549956 73788
rect 547880 33788 547932 33794
rect 547880 33730 547932 33736
rect 547892 16574 547920 33730
rect 545224 16546 545344 16574
rect 546512 16546 547552 16574
rect 547892 16546 548656 16574
rect 545120 1284 545172 1290
rect 545120 1226 545172 1232
rect 545316 480 545344 16546
rect 546408 1284 546460 1290
rect 546408 1226 546460 1232
rect 546420 480 546448 1226
rect 547524 480 547552 16546
rect 548628 480 548656 16546
rect 549720 15904 549772 15910
rect 549720 15846 549772 15852
rect 549732 480 549760 15846
rect 549916 3534 549944 73782
rect 553400 72480 553452 72486
rect 553400 72422 553452 72428
rect 552664 60036 552716 60042
rect 552664 59978 552716 59984
rect 552020 43444 552072 43450
rect 552020 43386 552072 43392
rect 552032 16574 552060 43386
rect 552032 16546 552612 16574
rect 550732 13116 550784 13122
rect 550732 13058 550784 13064
rect 549904 3528 549956 3534
rect 549904 3470 549956 3476
rect 550744 3398 550772 13058
rect 550824 3528 550876 3534
rect 550824 3470 550876 3476
rect 552584 3482 552612 16546
rect 552676 3670 552704 59978
rect 553412 16574 553440 72422
rect 553412 16546 554176 16574
rect 552664 3664 552716 3670
rect 552664 3606 552716 3612
rect 550732 3392 550784 3398
rect 550732 3334 550784 3340
rect 550836 480 550864 3470
rect 552584 3454 553072 3482
rect 551928 3392 551980 3398
rect 551928 3334 551980 3340
rect 551940 480 551968 3334
rect 553044 480 553072 3454
rect 554148 480 554176 16546
rect 555240 3664 555292 3670
rect 555240 3606 555292 3612
rect 555252 480 555280 3606
rect 556172 1290 556200 90306
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 88097 580212 88266
rect 580170 88088 580226 88097
rect 580170 88023 580226 88032
rect 580172 75880 580224 75886
rect 580172 75822 580224 75828
rect 580184 74905 580212 75822
rect 580170 74896 580226 74905
rect 580170 74831 580226 74840
rect 580172 62076 580224 62082
rect 580172 62018 580224 62024
rect 580184 61713 580212 62018
rect 580170 61704 580226 61713
rect 580170 61639 580226 61648
rect 580172 49700 580224 49706
rect 580172 49642 580224 49648
rect 580184 48521 580212 49642
rect 580170 48512 580226 48521
rect 580170 48447 580226 48456
rect 556252 42084 556304 42090
rect 556252 42026 556304 42032
rect 556264 16574 556292 42026
rect 580172 35896 580224 35902
rect 580172 35838 580224 35844
rect 580184 35329 580212 35838
rect 580170 35320 580226 35329
rect 580170 35255 580226 35264
rect 557540 32428 557592 32434
rect 557540 32370 557592 32376
rect 557552 16574 557580 32370
rect 580172 23452 580224 23458
rect 580172 23394 580224 23400
rect 580184 22137 580212 23394
rect 580170 22128 580226 22137
rect 580170 22063 580226 22072
rect 556264 16546 556384 16574
rect 557552 16546 558592 16574
rect 556160 1284 556212 1290
rect 556160 1226 556212 1232
rect 556356 480 556384 16546
rect 557448 1284 557500 1290
rect 557448 1226 557500 1232
rect 557460 480 557488 1226
rect 558564 480 558592 16546
rect 580172 9648 580224 9654
rect 580172 9590 580224 9596
rect 580184 8945 580212 9590
rect 580170 8936 580226 8945
rect 580170 8871 580226 8880
rect 559656 4820 559708 4826
rect 559656 4762 559708 4768
rect 559668 480 559696 4762
rect 562968 3596 563020 3602
rect 562968 3538 563020 3544
rect 561864 3460 561916 3466
rect 561864 3402 561916 3408
rect 561876 480 561904 3402
rect 562980 480 563008 3538
rect 564070 3360 564126 3369
rect 564070 3295 564126 3304
rect 564084 480 564112 3295
rect 291354 326 291884 354
rect 291354 -960 291466 326
rect 292458 -960 292570 480
rect 293562 -960 293674 480
rect 294666 -960 294778 480
rect 295770 -960 295882 480
rect 296874 -960 296986 480
rect 297978 -960 298090 480
rect 299082 -960 299194 480
rect 300186 -960 300298 480
rect 301290 -960 301402 480
rect 302394 -960 302506 480
rect 303498 -960 303610 480
rect 304602 -960 304714 480
rect 305706 -960 305818 480
rect 306810 -960 306922 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310122 -960 310234 480
rect 311226 -960 311338 480
rect 312330 -960 312442 480
rect 313434 -960 313546 480
rect 314538 -960 314650 480
rect 315642 -960 315754 480
rect 316746 -960 316858 480
rect 317850 -960 317962 480
rect 318954 -960 319066 480
rect 320058 -960 320170 480
rect 321162 -960 321274 480
rect 322266 -960 322378 480
rect 323370 -960 323482 480
rect 324474 -960 324586 480
rect 325578 -960 325690 480
rect 326682 -960 326794 480
rect 327786 -960 327898 480
rect 328890 -960 329002 480
rect 329994 -960 330106 480
rect 331098 -960 331210 480
rect 332202 -960 332314 480
rect 333306 -960 333418 480
rect 334410 -960 334522 480
rect 335514 -960 335626 480
rect 336618 -960 336730 480
rect 337722 -960 337834 480
rect 338826 -960 338938 480
rect 339930 -960 340042 480
rect 341034 -960 341146 480
rect 342138 -960 342250 480
rect 343242 -960 343354 480
rect 344346 -960 344458 480
rect 345450 -960 345562 480
rect 346554 -960 346666 480
rect 347658 -960 347770 480
rect 348762 -960 348874 480
rect 349866 -960 349978 480
rect 350970 -960 351082 480
rect 352074 -960 352186 480
rect 353178 -960 353290 480
rect 354282 -960 354394 480
rect 355386 -960 355498 480
rect 356490 -960 356602 480
rect 357594 -960 357706 480
rect 358698 -960 358810 480
rect 359802 -960 359914 480
rect 360906 -960 361018 480
rect 362010 -960 362122 480
rect 363114 -960 363226 480
rect 364218 -960 364330 480
rect 365322 -960 365434 480
rect 366426 -960 366538 480
rect 367530 -960 367642 480
rect 368634 -960 368746 480
rect 369738 -960 369850 480
rect 370842 -960 370954 480
rect 371946 -960 372058 480
rect 373050 -960 373162 480
rect 374154 -960 374266 480
rect 375258 -960 375370 480
rect 376362 -960 376474 480
rect 377466 -960 377578 480
rect 378570 -960 378682 480
rect 379674 -960 379786 480
rect 380778 -960 380890 480
rect 381882 -960 381994 480
rect 382986 -960 383098 480
rect 384090 -960 384202 480
rect 385194 -960 385306 480
rect 386298 -960 386410 480
rect 387402 -960 387514 480
rect 388506 -960 388618 480
rect 389610 -960 389722 480
rect 390714 -960 390826 480
rect 391818 -960 391930 480
rect 392922 -960 393034 480
rect 394026 -960 394138 480
rect 395130 -960 395242 480
rect 396234 -960 396346 480
rect 397338 -960 397450 480
rect 398442 -960 398554 480
rect 399546 -960 399658 480
rect 400650 -960 400762 480
rect 401754 -960 401866 480
rect 402858 -960 402970 480
rect 403962 -960 404074 480
rect 405066 -960 405178 480
rect 406170 -960 406282 480
rect 407274 -960 407386 480
rect 408378 -960 408490 480
rect 409482 -960 409594 480
rect 410586 -960 410698 480
rect 411690 -960 411802 480
rect 412794 -960 412906 480
rect 413898 -960 414010 480
rect 415002 -960 415114 480
rect 416106 -960 416218 480
rect 417210 -960 417322 480
rect 418314 -960 418426 480
rect 419418 -960 419530 480
rect 420522 -960 420634 480
rect 421626 -960 421738 480
rect 422730 -960 422842 480
rect 423834 -960 423946 480
rect 424938 -960 425050 480
rect 426042 -960 426154 480
rect 427146 -960 427258 480
rect 428250 -960 428362 480
rect 429354 -960 429466 480
rect 430458 -960 430570 480
rect 431562 -960 431674 480
rect 432666 -960 432778 480
rect 433770 -960 433882 480
rect 434874 -960 434986 480
rect 435978 -960 436090 480
rect 437082 -960 437194 480
rect 438186 -960 438298 480
rect 439290 -960 439402 480
rect 440394 -960 440506 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443706 -960 443818 480
rect 444810 -960 444922 480
rect 445914 -960 446026 480
rect 447018 -960 447130 480
rect 448122 -960 448234 480
rect 449226 -960 449338 480
rect 450330 -960 450442 480
rect 451434 -960 451546 480
rect 452538 -960 452650 480
rect 453642 -960 453754 480
rect 454746 -960 454858 480
rect 455850 -960 455962 480
rect 456954 -960 457066 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460266 -960 460378 480
rect 461370 -960 461482 480
rect 462474 -960 462586 480
rect 463578 -960 463690 480
rect 464682 -960 464794 480
rect 465786 -960 465898 480
rect 466890 -960 467002 480
rect 467994 -960 468106 480
rect 469098 -960 469210 480
rect 470202 -960 470314 480
rect 471306 -960 471418 480
rect 472410 -960 472522 480
rect 473514 -960 473626 480
rect 474618 -960 474730 480
rect 475722 -960 475834 480
rect 476826 -960 476938 480
rect 477930 -960 478042 480
rect 479034 -960 479146 480
rect 480138 -960 480250 480
rect 481242 -960 481354 480
rect 482346 -960 482458 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485658 -960 485770 480
rect 486762 -960 486874 480
rect 487866 -960 487978 480
rect 488970 -960 489082 480
rect 490074 -960 490186 480
rect 491178 -960 491290 480
rect 492282 -960 492394 480
rect 493386 -960 493498 480
rect 494490 -960 494602 480
rect 495594 -960 495706 480
rect 496698 -960 496810 480
rect 497802 -960 497914 480
rect 498906 -960 499018 480
rect 500010 -960 500122 480
rect 501114 -960 501226 480
rect 502218 -960 502330 480
rect 503322 -960 503434 480
rect 504426 -960 504538 480
rect 505530 -960 505642 480
rect 506634 -960 506746 480
rect 507738 -960 507850 480
rect 508842 -960 508954 480
rect 509946 -960 510058 480
rect 511050 -960 511162 480
rect 512154 -960 512266 480
rect 513258 -960 513370 480
rect 514362 -960 514474 480
rect 515466 -960 515578 480
rect 516570 -960 516682 480
rect 517674 -960 517786 480
rect 518778 -960 518890 480
rect 519882 -960 519994 480
rect 520986 -960 521098 480
rect 522090 -960 522202 480
rect 523194 -960 523306 480
rect 524298 -960 524410 480
rect 525402 -960 525514 480
rect 526506 -960 526618 480
rect 527610 -960 527722 480
rect 528714 -960 528826 480
rect 529818 -960 529930 480
rect 530922 -960 531034 480
rect 532026 -960 532138 480
rect 533130 -960 533242 480
rect 534234 -960 534346 480
rect 535338 -960 535450 480
rect 536442 -960 536554 480
rect 537546 -960 537658 480
rect 538650 -960 538762 480
rect 539754 -960 539866 480
rect 540858 -960 540970 480
rect 541962 -960 542074 480
rect 543066 -960 543178 480
rect 544170 -960 544282 480
rect 545274 -960 545386 480
rect 546378 -960 546490 480
rect 547482 -960 547594 480
rect 548586 -960 548698 480
rect 549690 -960 549802 480
rect 550794 -960 550906 480
rect 551898 -960 552010 480
rect 553002 -960 553114 480
rect 554106 -960 554218 480
rect 555210 -960 555322 480
rect 556314 -960 556426 480
rect 557418 -960 557530 480
rect 558522 -960 558634 480
rect 559626 -960 559738 480
rect 560730 -960 560842 480
rect 561834 -960 561946 480
rect 562938 -960 563050 480
rect 564042 -960 564154 480
<< via2 >>
rect 2778 681400 2834 681456
rect 3422 668480 3478 668536
rect 3330 616800 3386 616856
rect 3330 603880 3386 603936
rect 3330 578040 3386 578096
rect 3330 526360 3386 526416
rect 3330 513440 3386 513496
rect 2962 500520 3018 500576
rect 3238 474680 3294 474736
rect 2962 423000 3018 423056
rect 3330 410080 3386 410136
rect 2962 397160 3018 397216
rect 3330 371320 3386 371376
rect 3330 319640 3386 319696
rect 3330 306720 3386 306776
rect 3330 293800 3386 293856
rect 3330 267960 3386 268016
rect 3514 655560 3570 655616
rect 3330 255040 3386 255096
rect 3606 629720 3662 629776
rect 3606 565120 3662 565176
rect 3422 242120 3478 242176
rect 3698 552200 3754 552256
rect 3790 461760 3846 461816
rect 3514 216280 3570 216336
rect 3882 448840 3938 448896
rect 3974 358400 4030 358456
rect 3606 203360 3662 203416
rect 3698 190440 3754 190496
rect 3422 151680 3478 151736
rect 4066 345480 4122 345536
rect 580262 694864 580318 694920
rect 580170 681672 580226 681728
rect 230386 257896 230442 257952
rect 353298 257624 353354 257680
rect 580170 668480 580226 668536
rect 230386 254088 230442 254144
rect 353942 254088 353998 254144
rect 353298 250552 353354 250608
rect 230386 250280 230442 250336
rect 353298 247016 353354 247072
rect 229650 246472 229706 246528
rect 353298 243480 353354 243536
rect 229282 242664 229338 242720
rect 353298 239944 353354 240000
rect 230018 238856 230074 238912
rect 353298 236408 353354 236464
rect 230202 235048 230258 235104
rect 353298 232872 353354 232928
rect 230386 231240 230442 231296
rect 353298 229336 353354 229392
rect 230386 227432 230442 227488
rect 353298 225800 353354 225856
rect 229650 223624 229706 223680
rect 353298 222264 353354 222320
rect 230386 219816 230442 219872
rect 353298 218728 353354 218784
rect 230386 216008 230442 216064
rect 353298 215228 353300 215248
rect 353300 215228 353352 215248
rect 353352 215228 353354 215248
rect 353298 215192 353354 215228
rect 230386 212200 230442 212256
rect 353298 211656 353354 211712
rect 229650 208392 229706 208448
rect 353298 208156 353300 208176
rect 353300 208156 353352 208176
rect 353352 208156 353354 208176
rect 353298 208120 353354 208156
rect 229466 204584 229522 204640
rect 353298 204584 353354 204640
rect 353298 201048 353354 201104
rect 230386 200776 230442 200832
rect 353298 197512 353354 197568
rect 229834 196968 229890 197024
rect 353298 193976 353354 194032
rect 230386 193180 230442 193216
rect 230386 193160 230388 193180
rect 230388 193160 230440 193180
rect 230440 193160 230442 193180
rect 230386 189352 230442 189408
rect 353298 186904 353354 186960
rect 230386 185544 230442 185600
rect 353298 183368 353354 183424
rect 229834 181736 229890 181792
rect 353298 179832 353354 179888
rect 230386 177964 230388 177984
rect 230388 177964 230440 177984
rect 230440 177964 230442 177984
rect 230386 177928 230442 177964
rect 353298 176296 353354 176352
rect 230386 174120 230442 174176
rect 353298 172760 353354 172816
rect 230386 170312 230442 170368
rect 230386 166504 230442 166560
rect 353298 165688 353354 165744
rect 3790 164600 3846 164656
rect 230386 162696 230442 162752
rect 353298 162152 353354 162208
rect 230386 158888 230442 158944
rect 354034 190440 354090 190496
rect 353942 158616 353998 158672
rect 229282 155080 229338 155136
rect 353298 155080 353354 155136
rect 353298 151544 353354 151600
rect 230386 151272 230442 151328
rect 230386 147464 230442 147520
rect 353298 144472 353354 144528
rect 230018 143656 230074 143712
rect 579894 642096 579950 642152
rect 579894 628904 579950 628960
rect 580170 615712 580226 615768
rect 580170 562944 580226 563000
rect 580170 536560 580226 536616
rect 580170 523368 580226 523424
rect 579618 510176 579674 510232
rect 580170 457408 580226 457464
rect 579802 431024 579858 431080
rect 579618 417832 579674 417888
rect 580170 404640 580226 404696
rect 580170 365064 580226 365120
rect 580170 325488 580226 325544
rect 580170 312296 580226 312352
rect 579986 272720 580042 272776
rect 580170 259528 580226 259584
rect 580354 589328 580410 589384
rect 580262 246336 580318 246392
rect 580170 219952 580226 220008
rect 579618 180376 579674 180432
rect 354126 169224 354182 169280
rect 580446 576136 580502 576192
rect 580538 483792 580594 483848
rect 580354 233144 580410 233200
rect 580630 470600 580686 470656
rect 580722 378256 580778 378312
rect 580446 206760 580502 206816
rect 580814 351872 580870 351928
rect 580538 193568 580594 193624
rect 579618 153992 579674 154048
rect 580906 299104 580962 299160
rect 580630 167184 580686 167240
rect 354034 148008 354090 148064
rect 353942 140936 353998 140992
rect 580170 140820 580226 140856
rect 580170 140800 580172 140820
rect 580172 140800 580224 140820
rect 580224 140800 580226 140820
rect 230386 139848 230442 139904
rect 3422 138760 3478 138816
rect 353298 137400 353354 137456
rect 229650 136040 229706 136096
rect 354218 133864 354274 133920
rect 229742 132232 229798 132288
rect 3146 112920 3202 112976
rect 3330 87080 3386 87136
rect 3330 74160 3386 74216
rect 3238 48320 3294 48376
rect 3330 35400 3386 35456
rect 353942 130328 353998 130384
rect 230386 128424 230442 128480
rect 230110 124616 230166 124672
rect 230018 120808 230074 120864
rect 229926 113192 229982 113248
rect 229834 109384 229890 109440
rect 229742 101768 229798 101824
rect 3606 100000 3662 100056
rect 3514 61240 3570 61296
rect 3422 22480 3478 22536
rect 3422 9596 3424 9616
rect 3424 9596 3476 9616
rect 3476 9596 3478 9616
rect 3422 9560 3478 9596
rect 24214 3304 24270 3360
rect 230386 117000 230442 117056
rect 580170 127608 580226 127664
rect 354586 126792 354642 126848
rect 354494 123256 354550 123312
rect 354402 119720 354458 119776
rect 354310 116184 354366 116240
rect 354218 112648 354274 112704
rect 354126 109112 354182 109168
rect 230386 105576 230442 105632
rect 354034 105576 354090 105632
rect 353942 102040 353998 102096
rect 247498 3576 247554 3632
rect 337106 3576 337162 3632
rect 580170 114452 580172 114472
rect 580172 114452 580224 114472
rect 580224 114452 580226 114472
rect 580170 114416 580226 114452
rect 579986 101224 580042 101280
rect 580170 88032 580226 88088
rect 580170 74840 580226 74896
rect 580170 61648 580226 61704
rect 580170 48456 580226 48512
rect 580170 35264 580226 35320
rect 580170 22072 580226 22128
rect 580170 8880 580226 8936
rect 564070 3304 564126 3360
<< metal3 >>
rect 580257 694922 580323 694925
rect 583520 694922 584960 695012
rect 580257 694920 584960 694922
rect 580257 694864 580262 694920
rect 580318 694864 584960 694920
rect 580257 694862 584960 694864
rect 580257 694859 580323 694862
rect 583520 694772 584960 694862
rect -960 694228 480 694468
rect 580165 681730 580231 681733
rect 583520 681730 584960 681820
rect 580165 681728 584960 681730
rect 580165 681672 580170 681728
rect 580226 681672 584960 681728
rect 580165 681670 584960 681672
rect 580165 681667 580231 681670
rect 583520 681580 584960 681670
rect -960 681458 480 681548
rect 2773 681458 2839 681461
rect -960 681456 2839 681458
rect -960 681400 2778 681456
rect 2834 681400 2839 681456
rect -960 681398 2839 681400
rect -960 681308 480 681398
rect 2773 681395 2839 681398
rect -960 668538 480 668628
rect 3417 668538 3483 668541
rect -960 668536 3483 668538
rect -960 668480 3422 668536
rect 3478 668480 3483 668536
rect -960 668478 3483 668480
rect -960 668388 480 668478
rect 3417 668475 3483 668478
rect 580165 668538 580231 668541
rect 583520 668538 584960 668628
rect 580165 668536 584960 668538
rect 580165 668480 580170 668536
rect 580226 668480 584960 668536
rect 580165 668478 584960 668480
rect 580165 668475 580231 668478
rect 583520 668388 584960 668478
rect -960 655618 480 655708
rect 3509 655618 3575 655621
rect -960 655616 3575 655618
rect -960 655560 3514 655616
rect 3570 655560 3575 655616
rect -960 655558 3575 655560
rect -960 655468 480 655558
rect 3509 655555 3575 655558
rect 583520 655196 584960 655436
rect -960 642548 480 642788
rect 579889 642154 579955 642157
rect 583520 642154 584960 642244
rect 579889 642152 584960 642154
rect 579889 642096 579894 642152
rect 579950 642096 584960 642152
rect 579889 642094 584960 642096
rect 579889 642091 579955 642094
rect 583520 642004 584960 642094
rect -960 629778 480 629868
rect 3601 629778 3667 629781
rect -960 629776 3667 629778
rect -960 629720 3606 629776
rect 3662 629720 3667 629776
rect -960 629718 3667 629720
rect -960 629628 480 629718
rect 3601 629715 3667 629718
rect 579889 628962 579955 628965
rect 583520 628962 584960 629052
rect 579889 628960 584960 628962
rect 579889 628904 579894 628960
rect 579950 628904 584960 628960
rect 579889 628902 584960 628904
rect 579889 628899 579955 628902
rect 583520 628812 584960 628902
rect -960 616858 480 616948
rect 3325 616858 3391 616861
rect -960 616856 3391 616858
rect -960 616800 3330 616856
rect 3386 616800 3391 616856
rect -960 616798 3391 616800
rect -960 616708 480 616798
rect 3325 616795 3391 616798
rect 580165 615770 580231 615773
rect 583520 615770 584960 615860
rect 580165 615768 584960 615770
rect 580165 615712 580170 615768
rect 580226 615712 584960 615768
rect 580165 615710 584960 615712
rect 580165 615707 580231 615710
rect 583520 615620 584960 615710
rect -960 603938 480 604028
rect 3325 603938 3391 603941
rect -960 603936 3391 603938
rect -960 603880 3330 603936
rect 3386 603880 3391 603936
rect -960 603878 3391 603880
rect -960 603788 480 603878
rect 3325 603875 3391 603878
rect 583520 602428 584960 602668
rect -960 590868 480 591108
rect 580349 589386 580415 589389
rect 583520 589386 584960 589476
rect 580349 589384 584960 589386
rect 580349 589328 580354 589384
rect 580410 589328 584960 589384
rect 580349 589326 584960 589328
rect 580349 589323 580415 589326
rect 583520 589236 584960 589326
rect -960 578098 480 578188
rect 3325 578098 3391 578101
rect -960 578096 3391 578098
rect -960 578040 3330 578096
rect 3386 578040 3391 578096
rect -960 578038 3391 578040
rect -960 577948 480 578038
rect 3325 578035 3391 578038
rect 580441 576194 580507 576197
rect 583520 576194 584960 576284
rect 580441 576192 584960 576194
rect 580441 576136 580446 576192
rect 580502 576136 584960 576192
rect 580441 576134 584960 576136
rect 580441 576131 580507 576134
rect 583520 576044 584960 576134
rect -960 565178 480 565268
rect 3601 565178 3667 565181
rect -960 565176 3667 565178
rect -960 565120 3606 565176
rect 3662 565120 3667 565176
rect -960 565118 3667 565120
rect -960 565028 480 565118
rect 3601 565115 3667 565118
rect 580165 563002 580231 563005
rect 583520 563002 584960 563092
rect 580165 563000 584960 563002
rect 580165 562944 580170 563000
rect 580226 562944 584960 563000
rect 580165 562942 584960 562944
rect 580165 562939 580231 562942
rect 583520 562852 584960 562942
rect -960 552258 480 552348
rect 3693 552258 3759 552261
rect -960 552256 3759 552258
rect -960 552200 3698 552256
rect 3754 552200 3759 552256
rect -960 552198 3759 552200
rect -960 552108 480 552198
rect 3693 552195 3759 552198
rect 583520 549660 584960 549900
rect -960 539188 480 539428
rect 580165 536618 580231 536621
rect 583520 536618 584960 536708
rect 580165 536616 584960 536618
rect 580165 536560 580170 536616
rect 580226 536560 584960 536616
rect 580165 536558 584960 536560
rect 580165 536555 580231 536558
rect 583520 536468 584960 536558
rect -960 526418 480 526508
rect 3325 526418 3391 526421
rect -960 526416 3391 526418
rect -960 526360 3330 526416
rect 3386 526360 3391 526416
rect -960 526358 3391 526360
rect -960 526268 480 526358
rect 3325 526355 3391 526358
rect 580165 523426 580231 523429
rect 583520 523426 584960 523516
rect 580165 523424 584960 523426
rect 580165 523368 580170 523424
rect 580226 523368 584960 523424
rect 580165 523366 584960 523368
rect 580165 523363 580231 523366
rect 583520 523276 584960 523366
rect -960 513498 480 513588
rect 3325 513498 3391 513501
rect -960 513496 3391 513498
rect -960 513440 3330 513496
rect 3386 513440 3391 513496
rect -960 513438 3391 513440
rect -960 513348 480 513438
rect 3325 513435 3391 513438
rect 579613 510234 579679 510237
rect 583520 510234 584960 510324
rect 579613 510232 584960 510234
rect 579613 510176 579618 510232
rect 579674 510176 584960 510232
rect 579613 510174 584960 510176
rect 579613 510171 579679 510174
rect 583520 510084 584960 510174
rect -960 500578 480 500668
rect 2957 500578 3023 500581
rect -960 500576 3023 500578
rect -960 500520 2962 500576
rect 3018 500520 3023 500576
rect -960 500518 3023 500520
rect -960 500428 480 500518
rect 2957 500515 3023 500518
rect 583520 496892 584960 497132
rect -960 487508 480 487748
rect 580533 483850 580599 483853
rect 583520 483850 584960 483940
rect 580533 483848 584960 483850
rect 580533 483792 580538 483848
rect 580594 483792 584960 483848
rect 580533 483790 584960 483792
rect 580533 483787 580599 483790
rect 583520 483700 584960 483790
rect -960 474738 480 474828
rect 3233 474738 3299 474741
rect -960 474736 3299 474738
rect -960 474680 3238 474736
rect 3294 474680 3299 474736
rect -960 474678 3299 474680
rect -960 474588 480 474678
rect 3233 474675 3299 474678
rect 580625 470658 580691 470661
rect 583520 470658 584960 470748
rect 580625 470656 584960 470658
rect 580625 470600 580630 470656
rect 580686 470600 584960 470656
rect 580625 470598 584960 470600
rect 580625 470595 580691 470598
rect 583520 470508 584960 470598
rect -960 461818 480 461908
rect 3785 461818 3851 461821
rect -960 461816 3851 461818
rect -960 461760 3790 461816
rect 3846 461760 3851 461816
rect -960 461758 3851 461760
rect -960 461668 480 461758
rect 3785 461755 3851 461758
rect 580165 457466 580231 457469
rect 583520 457466 584960 457556
rect 580165 457464 584960 457466
rect 580165 457408 580170 457464
rect 580226 457408 584960 457464
rect 580165 457406 584960 457408
rect 580165 457403 580231 457406
rect 583520 457316 584960 457406
rect -960 448898 480 448988
rect 3877 448898 3943 448901
rect -960 448896 3943 448898
rect -960 448840 3882 448896
rect 3938 448840 3943 448896
rect -960 448838 3943 448840
rect -960 448748 480 448838
rect 3877 448835 3943 448838
rect 583520 444124 584960 444364
rect -960 435828 480 436068
rect 579797 431082 579863 431085
rect 583520 431082 584960 431172
rect 579797 431080 584960 431082
rect 579797 431024 579802 431080
rect 579858 431024 584960 431080
rect 579797 431022 584960 431024
rect 579797 431019 579863 431022
rect 583520 430932 584960 431022
rect -960 423058 480 423148
rect 2957 423058 3023 423061
rect -960 423056 3023 423058
rect -960 423000 2962 423056
rect 3018 423000 3023 423056
rect -960 422998 3023 423000
rect -960 422908 480 422998
rect 2957 422995 3023 422998
rect 579613 417890 579679 417893
rect 583520 417890 584960 417980
rect 579613 417888 584960 417890
rect 579613 417832 579618 417888
rect 579674 417832 584960 417888
rect 579613 417830 584960 417832
rect 579613 417827 579679 417830
rect 583520 417740 584960 417830
rect -960 410138 480 410228
rect 3325 410138 3391 410141
rect -960 410136 3391 410138
rect -960 410080 3330 410136
rect 3386 410080 3391 410136
rect -960 410078 3391 410080
rect -960 409988 480 410078
rect 3325 410075 3391 410078
rect 580165 404698 580231 404701
rect 583520 404698 584960 404788
rect 580165 404696 584960 404698
rect 580165 404640 580170 404696
rect 580226 404640 584960 404696
rect 580165 404638 584960 404640
rect 580165 404635 580231 404638
rect 583520 404548 584960 404638
rect -960 397218 480 397308
rect 2957 397218 3023 397221
rect -960 397216 3023 397218
rect -960 397160 2962 397216
rect 3018 397160 3023 397216
rect -960 397158 3023 397160
rect -960 397068 480 397158
rect 2957 397155 3023 397158
rect 583520 391356 584960 391596
rect -960 384148 480 384388
rect 580717 378314 580783 378317
rect 583520 378314 584960 378404
rect 580717 378312 584960 378314
rect 580717 378256 580722 378312
rect 580778 378256 584960 378312
rect 580717 378254 584960 378256
rect 580717 378251 580783 378254
rect 583520 378164 584960 378254
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3969 358458 4035 358461
rect -960 358456 4035 358458
rect -960 358400 3974 358456
rect 4030 358400 4035 358456
rect -960 358398 4035 358400
rect -960 358308 480 358398
rect 3969 358395 4035 358398
rect 580809 351930 580875 351933
rect 583520 351930 584960 352020
rect 580809 351928 584960 351930
rect 580809 351872 580814 351928
rect 580870 351872 584960 351928
rect 580809 351870 584960 351872
rect 580809 351867 580875 351870
rect 583520 351780 584960 351870
rect -960 345538 480 345628
rect 4061 345538 4127 345541
rect -960 345536 4127 345538
rect -960 345480 4066 345536
rect 4122 345480 4127 345536
rect -960 345478 4127 345480
rect -960 345388 480 345478
rect 4061 345475 4127 345478
rect 583520 338588 584960 338828
rect -960 332468 480 332708
rect 580165 325546 580231 325549
rect 583520 325546 584960 325636
rect 580165 325544 584960 325546
rect 580165 325488 580170 325544
rect 580226 325488 584960 325544
rect 580165 325486 584960 325488
rect 580165 325483 580231 325486
rect 583520 325396 584960 325486
rect -960 319698 480 319788
rect 3325 319698 3391 319701
rect -960 319696 3391 319698
rect -960 319640 3330 319696
rect 3386 319640 3391 319696
rect -960 319638 3391 319640
rect -960 319548 480 319638
rect 3325 319635 3391 319638
rect 580165 312354 580231 312357
rect 583520 312354 584960 312444
rect 580165 312352 584960 312354
rect 580165 312296 580170 312352
rect 580226 312296 584960 312352
rect 580165 312294 584960 312296
rect 580165 312291 580231 312294
rect 583520 312204 584960 312294
rect -960 306778 480 306868
rect 3325 306778 3391 306781
rect -960 306776 3391 306778
rect -960 306720 3330 306776
rect 3386 306720 3391 306776
rect -960 306718 3391 306720
rect -960 306628 480 306718
rect 3325 306715 3391 306718
rect 580901 299162 580967 299165
rect 583520 299162 584960 299252
rect 580901 299160 584960 299162
rect 580901 299104 580906 299160
rect 580962 299104 584960 299160
rect 580901 299102 584960 299104
rect 580901 299099 580967 299102
rect 583520 299012 584960 299102
rect -960 293858 480 293948
rect 3325 293858 3391 293861
rect -960 293856 3391 293858
rect -960 293800 3330 293856
rect 3386 293800 3391 293856
rect -960 293798 3391 293800
rect -960 293708 480 293798
rect 3325 293795 3391 293798
rect 583520 285820 584960 286060
rect -960 280788 480 281028
rect 579981 272778 580047 272781
rect 583520 272778 584960 272868
rect 579981 272776 584960 272778
rect 579981 272720 579986 272776
rect 580042 272720 584960 272776
rect 579981 272718 584960 272720
rect 579981 272715 580047 272718
rect 583520 272628 584960 272718
rect -960 268018 480 268108
rect 3325 268018 3391 268021
rect -960 268016 3391 268018
rect -960 267960 3330 268016
rect 3386 267960 3391 268016
rect -960 267958 3391 267960
rect -960 267868 480 267958
rect 3325 267955 3391 267958
rect 580165 259586 580231 259589
rect 583520 259586 584960 259676
rect 580165 259584 584960 259586
rect 580165 259528 580170 259584
rect 580226 259528 584960 259584
rect 580165 259526 584960 259528
rect 580165 259523 580231 259526
rect 583520 259436 584960 259526
rect 230381 257954 230447 257957
rect 230381 257952 232116 257954
rect 230381 257896 230386 257952
rect 230442 257896 232116 257952
rect 230381 257894 232116 257896
rect 230381 257891 230447 257894
rect 353293 257682 353359 257685
rect 351900 257680 353359 257682
rect 351900 257624 353298 257680
rect 353354 257624 353359 257680
rect 351900 257622 353359 257624
rect 353293 257619 353359 257622
rect -960 255098 480 255188
rect 3325 255098 3391 255101
rect -960 255096 3391 255098
rect -960 255040 3330 255096
rect 3386 255040 3391 255096
rect -960 255038 3391 255040
rect -960 254948 480 255038
rect 3325 255035 3391 255038
rect 230381 254146 230447 254149
rect 353937 254146 354003 254149
rect 230381 254144 232116 254146
rect 230381 254088 230386 254144
rect 230442 254088 232116 254144
rect 230381 254086 232116 254088
rect 351900 254144 354003 254146
rect 351900 254088 353942 254144
rect 353998 254088 354003 254144
rect 351900 254086 354003 254088
rect 230381 254083 230447 254086
rect 353937 254083 354003 254086
rect 353293 250610 353359 250613
rect 351900 250608 353359 250610
rect 351900 250552 353298 250608
rect 353354 250552 353359 250608
rect 351900 250550 353359 250552
rect 353293 250547 353359 250550
rect 230381 250338 230447 250341
rect 230381 250336 232116 250338
rect 230381 250280 230386 250336
rect 230442 250280 232116 250336
rect 230381 250278 232116 250280
rect 230381 250275 230447 250278
rect 353293 247074 353359 247077
rect 351900 247072 353359 247074
rect 351900 247016 353298 247072
rect 353354 247016 353359 247072
rect 351900 247014 353359 247016
rect 353293 247011 353359 247014
rect 229645 246530 229711 246533
rect 229645 246528 232116 246530
rect 229645 246472 229650 246528
rect 229706 246472 232116 246528
rect 229645 246470 232116 246472
rect 229645 246467 229711 246470
rect 580257 246394 580323 246397
rect 583520 246394 584960 246484
rect 580257 246392 584960 246394
rect 580257 246336 580262 246392
rect 580318 246336 584960 246392
rect 580257 246334 584960 246336
rect 580257 246331 580323 246334
rect 583520 246244 584960 246334
rect 353293 243538 353359 243541
rect 351900 243536 353359 243538
rect 351900 243480 353298 243536
rect 353354 243480 353359 243536
rect 351900 243478 353359 243480
rect 353293 243475 353359 243478
rect 229277 242722 229343 242725
rect 229277 242720 232116 242722
rect 229277 242664 229282 242720
rect 229338 242664 232116 242720
rect 229277 242662 232116 242664
rect 229277 242659 229343 242662
rect -960 242178 480 242268
rect 3417 242178 3483 242181
rect -960 242176 3483 242178
rect -960 242120 3422 242176
rect 3478 242120 3483 242176
rect -960 242118 3483 242120
rect -960 242028 480 242118
rect 3417 242115 3483 242118
rect 353293 240002 353359 240005
rect 351900 240000 353359 240002
rect 351900 239944 353298 240000
rect 353354 239944 353359 240000
rect 351900 239942 353359 239944
rect 353293 239939 353359 239942
rect 230013 238914 230079 238917
rect 230013 238912 232116 238914
rect 230013 238856 230018 238912
rect 230074 238856 232116 238912
rect 230013 238854 232116 238856
rect 230013 238851 230079 238854
rect 353293 236466 353359 236469
rect 351900 236464 353359 236466
rect 351900 236408 353298 236464
rect 353354 236408 353359 236464
rect 351900 236406 353359 236408
rect 353293 236403 353359 236406
rect 230197 235106 230263 235109
rect 230197 235104 232116 235106
rect 230197 235048 230202 235104
rect 230258 235048 232116 235104
rect 230197 235046 232116 235048
rect 230197 235043 230263 235046
rect 580349 233202 580415 233205
rect 583520 233202 584960 233292
rect 580349 233200 584960 233202
rect 580349 233144 580354 233200
rect 580410 233144 584960 233200
rect 580349 233142 584960 233144
rect 580349 233139 580415 233142
rect 583520 233052 584960 233142
rect 353293 232930 353359 232933
rect 351900 232928 353359 232930
rect 351900 232872 353298 232928
rect 353354 232872 353359 232928
rect 351900 232870 353359 232872
rect 353293 232867 353359 232870
rect 230381 231298 230447 231301
rect 230381 231296 232116 231298
rect 230381 231240 230386 231296
rect 230442 231240 232116 231296
rect 230381 231238 232116 231240
rect 230381 231235 230447 231238
rect 353293 229394 353359 229397
rect 351900 229392 353359 229394
rect -960 229108 480 229348
rect 351900 229336 353298 229392
rect 353354 229336 353359 229392
rect 351900 229334 353359 229336
rect 353293 229331 353359 229334
rect 230381 227490 230447 227493
rect 230381 227488 232116 227490
rect 230381 227432 230386 227488
rect 230442 227432 232116 227488
rect 230381 227430 232116 227432
rect 230381 227427 230447 227430
rect 353293 225858 353359 225861
rect 351900 225856 353359 225858
rect 351900 225800 353298 225856
rect 353354 225800 353359 225856
rect 351900 225798 353359 225800
rect 353293 225795 353359 225798
rect 229645 223682 229711 223685
rect 229645 223680 232116 223682
rect 229645 223624 229650 223680
rect 229706 223624 232116 223680
rect 229645 223622 232116 223624
rect 229645 223619 229711 223622
rect 353293 222322 353359 222325
rect 351900 222320 353359 222322
rect 351900 222264 353298 222320
rect 353354 222264 353359 222320
rect 351900 222262 353359 222264
rect 353293 222259 353359 222262
rect 580165 220010 580231 220013
rect 583520 220010 584960 220100
rect 580165 220008 584960 220010
rect 580165 219952 580170 220008
rect 580226 219952 584960 220008
rect 580165 219950 584960 219952
rect 580165 219947 580231 219950
rect 230381 219874 230447 219877
rect 230381 219872 232116 219874
rect 230381 219816 230386 219872
rect 230442 219816 232116 219872
rect 583520 219860 584960 219950
rect 230381 219814 232116 219816
rect 230381 219811 230447 219814
rect 353293 218786 353359 218789
rect 351900 218784 353359 218786
rect 351900 218728 353298 218784
rect 353354 218728 353359 218784
rect 351900 218726 353359 218728
rect 353293 218723 353359 218726
rect -960 216338 480 216428
rect 3509 216338 3575 216341
rect -960 216336 3575 216338
rect -960 216280 3514 216336
rect 3570 216280 3575 216336
rect -960 216278 3575 216280
rect -960 216188 480 216278
rect 3509 216275 3575 216278
rect 230381 216066 230447 216069
rect 230381 216064 232116 216066
rect 230381 216008 230386 216064
rect 230442 216008 232116 216064
rect 230381 216006 232116 216008
rect 230381 216003 230447 216006
rect 353293 215250 353359 215253
rect 351900 215248 353359 215250
rect 351900 215192 353298 215248
rect 353354 215192 353359 215248
rect 351900 215190 353359 215192
rect 353293 215187 353359 215190
rect 230381 212258 230447 212261
rect 230381 212256 232116 212258
rect 230381 212200 230386 212256
rect 230442 212200 232116 212256
rect 230381 212198 232116 212200
rect 230381 212195 230447 212198
rect 353293 211714 353359 211717
rect 351900 211712 353359 211714
rect 351900 211656 353298 211712
rect 353354 211656 353359 211712
rect 351900 211654 353359 211656
rect 353293 211651 353359 211654
rect 229645 208450 229711 208453
rect 229645 208448 232116 208450
rect 229645 208392 229650 208448
rect 229706 208392 232116 208448
rect 229645 208390 232116 208392
rect 229645 208387 229711 208390
rect 353293 208178 353359 208181
rect 351900 208176 353359 208178
rect 351900 208120 353298 208176
rect 353354 208120 353359 208176
rect 351900 208118 353359 208120
rect 353293 208115 353359 208118
rect 580441 206818 580507 206821
rect 583520 206818 584960 206908
rect 580441 206816 584960 206818
rect 580441 206760 580446 206816
rect 580502 206760 584960 206816
rect 580441 206758 584960 206760
rect 580441 206755 580507 206758
rect 583520 206668 584960 206758
rect 229461 204642 229527 204645
rect 353293 204642 353359 204645
rect 229461 204640 232116 204642
rect 229461 204584 229466 204640
rect 229522 204584 232116 204640
rect 229461 204582 232116 204584
rect 351900 204640 353359 204642
rect 351900 204584 353298 204640
rect 353354 204584 353359 204640
rect 351900 204582 353359 204584
rect 229461 204579 229527 204582
rect 353293 204579 353359 204582
rect -960 203418 480 203508
rect 3601 203418 3667 203421
rect -960 203416 3667 203418
rect -960 203360 3606 203416
rect 3662 203360 3667 203416
rect -960 203358 3667 203360
rect -960 203268 480 203358
rect 3601 203355 3667 203358
rect 353293 201106 353359 201109
rect 351900 201104 353359 201106
rect 351900 201048 353298 201104
rect 353354 201048 353359 201104
rect 351900 201046 353359 201048
rect 353293 201043 353359 201046
rect 230381 200834 230447 200837
rect 230381 200832 232116 200834
rect 230381 200776 230386 200832
rect 230442 200776 232116 200832
rect 230381 200774 232116 200776
rect 230381 200771 230447 200774
rect 353293 197570 353359 197573
rect 351900 197568 353359 197570
rect 351900 197512 353298 197568
rect 353354 197512 353359 197568
rect 351900 197510 353359 197512
rect 353293 197507 353359 197510
rect 229829 197026 229895 197029
rect 229829 197024 232116 197026
rect 229829 196968 229834 197024
rect 229890 196968 232116 197024
rect 229829 196966 232116 196968
rect 229829 196963 229895 196966
rect 353293 194034 353359 194037
rect 351900 194032 353359 194034
rect 351900 193976 353298 194032
rect 353354 193976 353359 194032
rect 351900 193974 353359 193976
rect 353293 193971 353359 193974
rect 580533 193626 580599 193629
rect 583520 193626 584960 193716
rect 580533 193624 584960 193626
rect 580533 193568 580538 193624
rect 580594 193568 584960 193624
rect 580533 193566 584960 193568
rect 580533 193563 580599 193566
rect 583520 193476 584960 193566
rect 230381 193218 230447 193221
rect 230381 193216 232116 193218
rect 230381 193160 230386 193216
rect 230442 193160 232116 193216
rect 230381 193158 232116 193160
rect 230381 193155 230447 193158
rect -960 190498 480 190588
rect 3693 190498 3759 190501
rect 354029 190498 354095 190501
rect -960 190496 3759 190498
rect -960 190440 3698 190496
rect 3754 190440 3759 190496
rect -960 190438 3759 190440
rect 351900 190496 354095 190498
rect 351900 190440 354034 190496
rect 354090 190440 354095 190496
rect 351900 190438 354095 190440
rect -960 190348 480 190438
rect 3693 190435 3759 190438
rect 354029 190435 354095 190438
rect 230381 189410 230447 189413
rect 230381 189408 232116 189410
rect 230381 189352 230386 189408
rect 230442 189352 232116 189408
rect 230381 189350 232116 189352
rect 230381 189347 230447 189350
rect 353293 186962 353359 186965
rect 351900 186960 353359 186962
rect 351900 186904 353298 186960
rect 353354 186904 353359 186960
rect 351900 186902 353359 186904
rect 353293 186899 353359 186902
rect 230381 185602 230447 185605
rect 230381 185600 232116 185602
rect 230381 185544 230386 185600
rect 230442 185544 232116 185600
rect 230381 185542 232116 185544
rect 230381 185539 230447 185542
rect 353293 183426 353359 183429
rect 351900 183424 353359 183426
rect 351900 183368 353298 183424
rect 353354 183368 353359 183424
rect 351900 183366 353359 183368
rect 353293 183363 353359 183366
rect 229829 181794 229895 181797
rect 229829 181792 232116 181794
rect 229829 181736 229834 181792
rect 229890 181736 232116 181792
rect 229829 181734 232116 181736
rect 229829 181731 229895 181734
rect 579613 180434 579679 180437
rect 583520 180434 584960 180524
rect 579613 180432 584960 180434
rect 579613 180376 579618 180432
rect 579674 180376 584960 180432
rect 579613 180374 584960 180376
rect 579613 180371 579679 180374
rect 583520 180284 584960 180374
rect 353293 179890 353359 179893
rect 351900 179888 353359 179890
rect 351900 179832 353298 179888
rect 353354 179832 353359 179888
rect 351900 179830 353359 179832
rect 353293 179827 353359 179830
rect 230381 177986 230447 177989
rect 230381 177984 232116 177986
rect 230381 177928 230386 177984
rect 230442 177928 232116 177984
rect 230381 177926 232116 177928
rect 230381 177923 230447 177926
rect -960 177428 480 177668
rect 353293 176354 353359 176357
rect 351900 176352 353359 176354
rect 351900 176296 353298 176352
rect 353354 176296 353359 176352
rect 351900 176294 353359 176296
rect 353293 176291 353359 176294
rect 230381 174178 230447 174181
rect 230381 174176 232116 174178
rect 230381 174120 230386 174176
rect 230442 174120 232116 174176
rect 230381 174118 232116 174120
rect 230381 174115 230447 174118
rect 353293 172818 353359 172821
rect 351900 172816 353359 172818
rect 351900 172760 353298 172816
rect 353354 172760 353359 172816
rect 351900 172758 353359 172760
rect 353293 172755 353359 172758
rect 230381 170370 230447 170373
rect 230381 170368 232116 170370
rect 230381 170312 230386 170368
rect 230442 170312 232116 170368
rect 230381 170310 232116 170312
rect 230381 170307 230447 170310
rect 354121 169282 354187 169285
rect 351900 169280 354187 169282
rect 351900 169224 354126 169280
rect 354182 169224 354187 169280
rect 351900 169222 354187 169224
rect 354121 169219 354187 169222
rect 580625 167242 580691 167245
rect 583520 167242 584960 167332
rect 580625 167240 584960 167242
rect 580625 167184 580630 167240
rect 580686 167184 584960 167240
rect 580625 167182 584960 167184
rect 580625 167179 580691 167182
rect 583520 167092 584960 167182
rect 230381 166562 230447 166565
rect 230381 166560 232116 166562
rect 230381 166504 230386 166560
rect 230442 166504 232116 166560
rect 230381 166502 232116 166504
rect 230381 166499 230447 166502
rect 353293 165746 353359 165749
rect 351900 165744 353359 165746
rect 351900 165688 353298 165744
rect 353354 165688 353359 165744
rect 351900 165686 353359 165688
rect 353293 165683 353359 165686
rect -960 164658 480 164748
rect 3785 164658 3851 164661
rect -960 164656 3851 164658
rect -960 164600 3790 164656
rect 3846 164600 3851 164656
rect -960 164598 3851 164600
rect -960 164508 480 164598
rect 3785 164595 3851 164598
rect 230381 162754 230447 162757
rect 230381 162752 232116 162754
rect 230381 162696 230386 162752
rect 230442 162696 232116 162752
rect 230381 162694 232116 162696
rect 230381 162691 230447 162694
rect 353293 162210 353359 162213
rect 351900 162208 353359 162210
rect 351900 162152 353298 162208
rect 353354 162152 353359 162208
rect 351900 162150 353359 162152
rect 353293 162147 353359 162150
rect 230381 158946 230447 158949
rect 230381 158944 232116 158946
rect 230381 158888 230386 158944
rect 230442 158888 232116 158944
rect 230381 158886 232116 158888
rect 230381 158883 230447 158886
rect 353937 158674 354003 158677
rect 351900 158672 354003 158674
rect 351900 158616 353942 158672
rect 353998 158616 354003 158672
rect 351900 158614 354003 158616
rect 353937 158611 354003 158614
rect 229277 155138 229343 155141
rect 353293 155138 353359 155141
rect 229277 155136 232116 155138
rect 229277 155080 229282 155136
rect 229338 155080 232116 155136
rect 229277 155078 232116 155080
rect 351900 155136 353359 155138
rect 351900 155080 353298 155136
rect 353354 155080 353359 155136
rect 351900 155078 353359 155080
rect 229277 155075 229343 155078
rect 353293 155075 353359 155078
rect 579613 154050 579679 154053
rect 583520 154050 584960 154140
rect 579613 154048 584960 154050
rect 579613 153992 579618 154048
rect 579674 153992 584960 154048
rect 579613 153990 584960 153992
rect 579613 153987 579679 153990
rect 583520 153900 584960 153990
rect -960 151738 480 151828
rect 3417 151738 3483 151741
rect -960 151736 3483 151738
rect -960 151680 3422 151736
rect 3478 151680 3483 151736
rect -960 151678 3483 151680
rect -960 151588 480 151678
rect 3417 151675 3483 151678
rect 353293 151602 353359 151605
rect 351900 151600 353359 151602
rect 351900 151544 353298 151600
rect 353354 151544 353359 151600
rect 351900 151542 353359 151544
rect 353293 151539 353359 151542
rect 230381 151330 230447 151333
rect 230381 151328 232116 151330
rect 230381 151272 230386 151328
rect 230442 151272 232116 151328
rect 230381 151270 232116 151272
rect 230381 151267 230447 151270
rect 354029 148066 354095 148069
rect 351900 148064 354095 148066
rect 351900 148008 354034 148064
rect 354090 148008 354095 148064
rect 351900 148006 354095 148008
rect 354029 148003 354095 148006
rect 230381 147522 230447 147525
rect 230381 147520 232116 147522
rect 230381 147464 230386 147520
rect 230442 147464 232116 147520
rect 230381 147462 232116 147464
rect 230381 147459 230447 147462
rect 353293 144530 353359 144533
rect 351900 144528 353359 144530
rect 351900 144472 353298 144528
rect 353354 144472 353359 144528
rect 351900 144470 353359 144472
rect 353293 144467 353359 144470
rect 230013 143714 230079 143717
rect 230013 143712 232116 143714
rect 230013 143656 230018 143712
rect 230074 143656 232116 143712
rect 230013 143654 232116 143656
rect 230013 143651 230079 143654
rect 353937 140994 354003 140997
rect 351900 140992 354003 140994
rect 351900 140936 353942 140992
rect 353998 140936 354003 140992
rect 351900 140934 354003 140936
rect 353937 140931 354003 140934
rect 580165 140858 580231 140861
rect 583520 140858 584960 140948
rect 580165 140856 584960 140858
rect 580165 140800 580170 140856
rect 580226 140800 584960 140856
rect 580165 140798 584960 140800
rect 580165 140795 580231 140798
rect 583520 140708 584960 140798
rect 230381 139906 230447 139909
rect 230381 139904 232116 139906
rect 230381 139848 230386 139904
rect 230442 139848 232116 139904
rect 230381 139846 232116 139848
rect 230381 139843 230447 139846
rect -960 138818 480 138908
rect 3417 138818 3483 138821
rect -960 138816 3483 138818
rect -960 138760 3422 138816
rect 3478 138760 3483 138816
rect -960 138758 3483 138760
rect -960 138668 480 138758
rect 3417 138755 3483 138758
rect 353293 137458 353359 137461
rect 351900 137456 353359 137458
rect 351900 137400 353298 137456
rect 353354 137400 353359 137456
rect 351900 137398 353359 137400
rect 353293 137395 353359 137398
rect 229645 136098 229711 136101
rect 229645 136096 232116 136098
rect 229645 136040 229650 136096
rect 229706 136040 232116 136096
rect 229645 136038 232116 136040
rect 229645 136035 229711 136038
rect 354213 133922 354279 133925
rect 351900 133920 354279 133922
rect 351900 133864 354218 133920
rect 354274 133864 354279 133920
rect 351900 133862 354279 133864
rect 354213 133859 354279 133862
rect 229737 132290 229803 132293
rect 229737 132288 232116 132290
rect 229737 132232 229742 132288
rect 229798 132232 232116 132288
rect 229737 132230 232116 132232
rect 229737 132227 229803 132230
rect 353937 130386 354003 130389
rect 351900 130384 354003 130386
rect 351900 130328 353942 130384
rect 353998 130328 354003 130384
rect 351900 130326 354003 130328
rect 353937 130323 354003 130326
rect 230381 128482 230447 128485
rect 230381 128480 232116 128482
rect 230381 128424 230386 128480
rect 230442 128424 232116 128480
rect 230381 128422 232116 128424
rect 230381 128419 230447 128422
rect 580165 127666 580231 127669
rect 583520 127666 584960 127756
rect 580165 127664 584960 127666
rect 580165 127608 580170 127664
rect 580226 127608 584960 127664
rect 580165 127606 584960 127608
rect 580165 127603 580231 127606
rect 583520 127516 584960 127606
rect 354581 126850 354647 126853
rect 351900 126848 354647 126850
rect 351900 126792 354586 126848
rect 354642 126792 354647 126848
rect 351900 126790 354647 126792
rect 354581 126787 354647 126790
rect -960 125748 480 125988
rect 230105 124674 230171 124677
rect 230105 124672 232116 124674
rect 230105 124616 230110 124672
rect 230166 124616 232116 124672
rect 230105 124614 232116 124616
rect 230105 124611 230171 124614
rect 354489 123314 354555 123317
rect 351900 123312 354555 123314
rect 351900 123256 354494 123312
rect 354550 123256 354555 123312
rect 351900 123254 354555 123256
rect 354489 123251 354555 123254
rect 230013 120866 230079 120869
rect 230013 120864 232116 120866
rect 230013 120808 230018 120864
rect 230074 120808 232116 120864
rect 230013 120806 232116 120808
rect 230013 120803 230079 120806
rect 354397 119778 354463 119781
rect 351900 119776 354463 119778
rect 351900 119720 354402 119776
rect 354458 119720 354463 119776
rect 351900 119718 354463 119720
rect 354397 119715 354463 119718
rect 230381 117058 230447 117061
rect 230381 117056 232116 117058
rect 230381 117000 230386 117056
rect 230442 117000 232116 117056
rect 230381 116998 232116 117000
rect 230381 116995 230447 116998
rect 354305 116242 354371 116245
rect 351900 116240 354371 116242
rect 351900 116184 354310 116240
rect 354366 116184 354371 116240
rect 351900 116182 354371 116184
rect 354305 116179 354371 116182
rect 580165 114474 580231 114477
rect 583520 114474 584960 114564
rect 580165 114472 584960 114474
rect 580165 114416 580170 114472
rect 580226 114416 584960 114472
rect 580165 114414 584960 114416
rect 580165 114411 580231 114414
rect 583520 114324 584960 114414
rect 229921 113250 229987 113253
rect 229921 113248 232116 113250
rect 229921 113192 229926 113248
rect 229982 113192 232116 113248
rect 229921 113190 232116 113192
rect 229921 113187 229987 113190
rect -960 112978 480 113068
rect 3141 112978 3207 112981
rect -960 112976 3207 112978
rect -960 112920 3146 112976
rect 3202 112920 3207 112976
rect -960 112918 3207 112920
rect -960 112828 480 112918
rect 3141 112915 3207 112918
rect 354213 112706 354279 112709
rect 351900 112704 354279 112706
rect 351900 112648 354218 112704
rect 354274 112648 354279 112704
rect 351900 112646 354279 112648
rect 354213 112643 354279 112646
rect 229829 109442 229895 109445
rect 229829 109440 232116 109442
rect 229829 109384 229834 109440
rect 229890 109384 232116 109440
rect 229829 109382 232116 109384
rect 229829 109379 229895 109382
rect 354121 109170 354187 109173
rect 351900 109168 354187 109170
rect 351900 109112 354126 109168
rect 354182 109112 354187 109168
rect 351900 109110 354187 109112
rect 354121 109107 354187 109110
rect 230381 105634 230447 105637
rect 354029 105634 354095 105637
rect 230381 105632 232116 105634
rect 230381 105576 230386 105632
rect 230442 105576 232116 105632
rect 230381 105574 232116 105576
rect 351900 105632 354095 105634
rect 351900 105576 354034 105632
rect 354090 105576 354095 105632
rect 351900 105574 354095 105576
rect 230381 105571 230447 105574
rect 354029 105571 354095 105574
rect 353937 102098 354003 102101
rect 351900 102096 354003 102098
rect 351900 102040 353942 102096
rect 353998 102040 354003 102096
rect 351900 102038 354003 102040
rect 353937 102035 354003 102038
rect 229737 101826 229803 101829
rect 229737 101824 232116 101826
rect 229737 101768 229742 101824
rect 229798 101768 232116 101824
rect 229737 101766 232116 101768
rect 229737 101763 229803 101766
rect 579981 101282 580047 101285
rect 583520 101282 584960 101372
rect 579981 101280 584960 101282
rect 579981 101224 579986 101280
rect 580042 101224 584960 101280
rect 579981 101222 584960 101224
rect 579981 101219 580047 101222
rect 583520 101132 584960 101222
rect -960 100058 480 100148
rect 3601 100058 3667 100061
rect -960 100056 3667 100058
rect -960 100000 3606 100056
rect 3662 100000 3667 100056
rect -960 99998 3667 100000
rect -960 99908 480 99998
rect 3601 99995 3667 99998
rect 580165 88090 580231 88093
rect 583520 88090 584960 88180
rect 580165 88088 584960 88090
rect 580165 88032 580170 88088
rect 580226 88032 584960 88088
rect 580165 88030 584960 88032
rect 580165 88027 580231 88030
rect 583520 87940 584960 88030
rect -960 87138 480 87228
rect 3325 87138 3391 87141
rect -960 87136 3391 87138
rect -960 87080 3330 87136
rect 3386 87080 3391 87136
rect -960 87078 3391 87080
rect -960 86988 480 87078
rect 3325 87075 3391 87078
rect 580165 74898 580231 74901
rect 583520 74898 584960 74988
rect 580165 74896 584960 74898
rect 580165 74840 580170 74896
rect 580226 74840 584960 74896
rect 580165 74838 584960 74840
rect 580165 74835 580231 74838
rect 583520 74748 584960 74838
rect -960 74218 480 74308
rect 3325 74218 3391 74221
rect -960 74216 3391 74218
rect -960 74160 3330 74216
rect 3386 74160 3391 74216
rect -960 74158 3391 74160
rect -960 74068 480 74158
rect 3325 74155 3391 74158
rect 580165 61706 580231 61709
rect 583520 61706 584960 61796
rect 580165 61704 584960 61706
rect 580165 61648 580170 61704
rect 580226 61648 584960 61704
rect 580165 61646 584960 61648
rect 580165 61643 580231 61646
rect 583520 61556 584960 61646
rect -960 61298 480 61388
rect 3509 61298 3575 61301
rect -960 61296 3575 61298
rect -960 61240 3514 61296
rect 3570 61240 3575 61296
rect -960 61238 3575 61240
rect -960 61148 480 61238
rect 3509 61235 3575 61238
rect 580165 48514 580231 48517
rect 583520 48514 584960 48604
rect 580165 48512 584960 48514
rect -960 48378 480 48468
rect 580165 48456 580170 48512
rect 580226 48456 584960 48512
rect 580165 48454 584960 48456
rect 580165 48451 580231 48454
rect 3233 48378 3299 48381
rect -960 48376 3299 48378
rect -960 48320 3238 48376
rect 3294 48320 3299 48376
rect 583520 48364 584960 48454
rect -960 48318 3299 48320
rect -960 48228 480 48318
rect 3233 48315 3299 48318
rect -960 35458 480 35548
rect 3325 35458 3391 35461
rect -960 35456 3391 35458
rect -960 35400 3330 35456
rect 3386 35400 3391 35456
rect -960 35398 3391 35400
rect -960 35308 480 35398
rect 3325 35395 3391 35398
rect 580165 35322 580231 35325
rect 583520 35322 584960 35412
rect 580165 35320 584960 35322
rect 580165 35264 580170 35320
rect 580226 35264 584960 35320
rect 580165 35262 584960 35264
rect 580165 35259 580231 35262
rect 583520 35172 584960 35262
rect -960 22538 480 22628
rect 3417 22538 3483 22541
rect -960 22536 3483 22538
rect -960 22480 3422 22536
rect 3478 22480 3483 22536
rect -960 22478 3483 22480
rect -960 22388 480 22478
rect 3417 22475 3483 22478
rect 580165 22130 580231 22133
rect 583520 22130 584960 22220
rect 580165 22128 584960 22130
rect 580165 22072 580170 22128
rect 580226 22072 584960 22128
rect 580165 22070 584960 22072
rect 580165 22067 580231 22070
rect 583520 21980 584960 22070
rect -960 9618 480 9708
rect 3417 9618 3483 9621
rect -960 9616 3483 9618
rect -960 9560 3422 9616
rect 3478 9560 3483 9616
rect -960 9558 3483 9560
rect -960 9468 480 9558
rect 3417 9555 3483 9558
rect 580165 8938 580231 8941
rect 583520 8938 584960 9028
rect 580165 8936 584960 8938
rect 580165 8880 580170 8936
rect 580226 8880 584960 8936
rect 580165 8878 584960 8880
rect 580165 8875 580231 8878
rect 583520 8788 584960 8878
rect 247493 3634 247559 3637
rect 238710 3632 247559 3634
rect 238710 3576 247498 3632
rect 247554 3576 247559 3632
rect 238710 3574 247559 3576
rect 24209 3362 24275 3365
rect 238710 3362 238770 3574
rect 247493 3571 247559 3574
rect 337101 3634 337167 3637
rect 337101 3632 345030 3634
rect 337101 3576 337106 3632
rect 337162 3576 345030 3632
rect 337101 3574 345030 3576
rect 337101 3571 337167 3574
rect 24209 3360 238770 3362
rect 24209 3304 24214 3360
rect 24270 3304 238770 3360
rect 24209 3302 238770 3304
rect 344970 3362 345030 3574
rect 564065 3362 564131 3365
rect 344970 3360 564131 3362
rect 344970 3304 564070 3360
rect 564126 3304 564131 3360
rect 344970 3302 564131 3304
rect 24209 3299 24275 3302
rect 564065 3299 564131 3302
<< metal4 >>
rect -9036 711868 -8416 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 -8416 711868
rect -9036 711548 -8416 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 -8416 711548
rect -9036 682954 -8416 711312
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 -8416 682954
rect -9036 682634 -8416 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 -8416 682634
rect -9036 646954 -8416 682398
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 -8416 646954
rect -9036 646634 -8416 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 -8416 646634
rect -9036 610954 -8416 646398
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 -8416 610954
rect -9036 610634 -8416 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 -8416 610634
rect -9036 574954 -8416 610398
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 -8416 574954
rect -9036 574634 -8416 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 -8416 574634
rect -9036 538954 -8416 574398
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 -8416 538954
rect -9036 538634 -8416 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 -8416 538634
rect -9036 502954 -8416 538398
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 -8416 502954
rect -9036 502634 -8416 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 -8416 502634
rect -9036 466954 -8416 502398
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 -8416 466954
rect -9036 466634 -8416 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 -8416 466634
rect -9036 430954 -8416 466398
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 -8416 430954
rect -9036 430634 -8416 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 -8416 430634
rect -9036 394954 -8416 430398
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 -8416 394954
rect -9036 394634 -8416 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 -8416 394634
rect -9036 358954 -8416 394398
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 -8416 358954
rect -9036 358634 -8416 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 -8416 358634
rect -9036 322954 -8416 358398
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 -8416 322954
rect -9036 322634 -8416 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 -8416 322634
rect -9036 286954 -8416 322398
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 -8416 286954
rect -9036 286634 -8416 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 -8416 286634
rect -9036 250954 -8416 286398
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 -8416 250954
rect -9036 250634 -8416 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 -8416 250634
rect -9036 214954 -8416 250398
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 -8416 214954
rect -9036 214634 -8416 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 -8416 214634
rect -9036 178954 -8416 214398
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 -8416 178954
rect -9036 178634 -8416 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 -8416 178634
rect -9036 142954 -8416 178398
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 -8416 142954
rect -9036 142634 -8416 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 -8416 142634
rect -9036 106954 -8416 142398
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 -8416 106954
rect -9036 106634 -8416 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 -8416 106634
rect -9036 70954 -8416 106398
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 -8416 70954
rect -9036 70634 -8416 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 -8416 70634
rect -9036 34954 -8416 70398
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 -8416 34954
rect -9036 34634 -8416 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 -8416 34634
rect -9036 -7376 -8416 34398
rect -8076 710908 -7456 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 -7456 710908
rect -8076 710588 -7456 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 -7456 710588
rect -8076 678454 -7456 710352
rect -8076 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 -7456 678454
rect -8076 678134 -7456 678218
rect -8076 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 -7456 678134
rect -8076 642454 -7456 677898
rect -8076 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 -7456 642454
rect -8076 642134 -7456 642218
rect -8076 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 -7456 642134
rect -8076 606454 -7456 641898
rect -8076 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 -7456 606454
rect -8076 606134 -7456 606218
rect -8076 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 -7456 606134
rect -8076 570454 -7456 605898
rect -8076 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 -7456 570454
rect -8076 570134 -7456 570218
rect -8076 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 -7456 570134
rect -8076 534454 -7456 569898
rect -8076 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 -7456 534454
rect -8076 534134 -7456 534218
rect -8076 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 -7456 534134
rect -8076 498454 -7456 533898
rect -8076 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 -7456 498454
rect -8076 498134 -7456 498218
rect -8076 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 -7456 498134
rect -8076 462454 -7456 497898
rect -8076 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 -7456 462454
rect -8076 462134 -7456 462218
rect -8076 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 -7456 462134
rect -8076 426454 -7456 461898
rect -8076 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 -7456 426454
rect -8076 426134 -7456 426218
rect -8076 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 -7456 426134
rect -8076 390454 -7456 425898
rect -8076 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 -7456 390454
rect -8076 390134 -7456 390218
rect -8076 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 -7456 390134
rect -8076 354454 -7456 389898
rect -8076 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 -7456 354454
rect -8076 354134 -7456 354218
rect -8076 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 -7456 354134
rect -8076 318454 -7456 353898
rect -8076 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 -7456 318454
rect -8076 318134 -7456 318218
rect -8076 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 -7456 318134
rect -8076 282454 -7456 317898
rect -8076 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 -7456 282454
rect -8076 282134 -7456 282218
rect -8076 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 -7456 282134
rect -8076 246454 -7456 281898
rect -8076 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 -7456 246454
rect -8076 246134 -7456 246218
rect -8076 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 -7456 246134
rect -8076 210454 -7456 245898
rect -8076 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 -7456 210454
rect -8076 210134 -7456 210218
rect -8076 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 -7456 210134
rect -8076 174454 -7456 209898
rect -8076 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 -7456 174454
rect -8076 174134 -7456 174218
rect -8076 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 -7456 174134
rect -8076 138454 -7456 173898
rect -8076 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 -7456 138454
rect -8076 138134 -7456 138218
rect -8076 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 -7456 138134
rect -8076 102454 -7456 137898
rect -8076 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 -7456 102454
rect -8076 102134 -7456 102218
rect -8076 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 -7456 102134
rect -8076 66454 -7456 101898
rect -8076 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 -7456 66454
rect -8076 66134 -7456 66218
rect -8076 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 -7456 66134
rect -8076 30454 -7456 65898
rect -8076 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 -7456 30454
rect -8076 30134 -7456 30218
rect -8076 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 -7456 30134
rect -8076 -6416 -7456 29898
rect -7116 709948 -6496 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 -6496 709948
rect -7116 709628 -6496 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 -6496 709628
rect -7116 673954 -6496 709392
rect -7116 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 -6496 673954
rect -7116 673634 -6496 673718
rect -7116 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 -6496 673634
rect -7116 637954 -6496 673398
rect -7116 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 -6496 637954
rect -7116 637634 -6496 637718
rect -7116 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 -6496 637634
rect -7116 601954 -6496 637398
rect -7116 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 -6496 601954
rect -7116 601634 -6496 601718
rect -7116 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 -6496 601634
rect -7116 565954 -6496 601398
rect -7116 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 -6496 565954
rect -7116 565634 -6496 565718
rect -7116 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 -6496 565634
rect -7116 529954 -6496 565398
rect -7116 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 -6496 529954
rect -7116 529634 -6496 529718
rect -7116 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 -6496 529634
rect -7116 493954 -6496 529398
rect -7116 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 -6496 493954
rect -7116 493634 -6496 493718
rect -7116 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 -6496 493634
rect -7116 457954 -6496 493398
rect -7116 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 -6496 457954
rect -7116 457634 -6496 457718
rect -7116 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 -6496 457634
rect -7116 421954 -6496 457398
rect -7116 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 -6496 421954
rect -7116 421634 -6496 421718
rect -7116 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 -6496 421634
rect -7116 385954 -6496 421398
rect -7116 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 -6496 385954
rect -7116 385634 -6496 385718
rect -7116 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 -6496 385634
rect -7116 349954 -6496 385398
rect -7116 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 -6496 349954
rect -7116 349634 -6496 349718
rect -7116 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 -6496 349634
rect -7116 313954 -6496 349398
rect -7116 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 -6496 313954
rect -7116 313634 -6496 313718
rect -7116 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 -6496 313634
rect -7116 277954 -6496 313398
rect -7116 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 -6496 277954
rect -7116 277634 -6496 277718
rect -7116 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 -6496 277634
rect -7116 241954 -6496 277398
rect -7116 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 -6496 241954
rect -7116 241634 -6496 241718
rect -7116 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 -6496 241634
rect -7116 205954 -6496 241398
rect -7116 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 -6496 205954
rect -7116 205634 -6496 205718
rect -7116 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 -6496 205634
rect -7116 169954 -6496 205398
rect -7116 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 -6496 169954
rect -7116 169634 -6496 169718
rect -7116 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 -6496 169634
rect -7116 133954 -6496 169398
rect -7116 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 -6496 133954
rect -7116 133634 -6496 133718
rect -7116 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 -6496 133634
rect -7116 97954 -6496 133398
rect -7116 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 -6496 97954
rect -7116 97634 -6496 97718
rect -7116 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 -6496 97634
rect -7116 61954 -6496 97398
rect -7116 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 -6496 61954
rect -7116 61634 -6496 61718
rect -7116 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 -6496 61634
rect -7116 25954 -6496 61398
rect -7116 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 -6496 25954
rect -7116 25634 -6496 25718
rect -7116 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 -6496 25634
rect -7116 -5456 -6496 25398
rect -6156 708988 -5536 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 -5536 708988
rect -6156 708668 -5536 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 -5536 708668
rect -6156 669454 -5536 708432
rect -6156 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 -5536 669454
rect -6156 669134 -5536 669218
rect -6156 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 -5536 669134
rect -6156 633454 -5536 668898
rect -6156 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 -5536 633454
rect -6156 633134 -5536 633218
rect -6156 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 -5536 633134
rect -6156 597454 -5536 632898
rect -6156 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 -5536 597454
rect -6156 597134 -5536 597218
rect -6156 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 -5536 597134
rect -6156 561454 -5536 596898
rect -6156 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 -5536 561454
rect -6156 561134 -5536 561218
rect -6156 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 -5536 561134
rect -6156 525454 -5536 560898
rect -6156 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 -5536 525454
rect -6156 525134 -5536 525218
rect -6156 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 -5536 525134
rect -6156 489454 -5536 524898
rect -6156 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 -5536 489454
rect -6156 489134 -5536 489218
rect -6156 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 -5536 489134
rect -6156 453454 -5536 488898
rect -6156 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 -5536 453454
rect -6156 453134 -5536 453218
rect -6156 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 -5536 453134
rect -6156 417454 -5536 452898
rect -6156 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 -5536 417454
rect -6156 417134 -5536 417218
rect -6156 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 -5536 417134
rect -6156 381454 -5536 416898
rect -6156 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 -5536 381454
rect -6156 381134 -5536 381218
rect -6156 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 -5536 381134
rect -6156 345454 -5536 380898
rect -6156 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 -5536 345454
rect -6156 345134 -5536 345218
rect -6156 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 -5536 345134
rect -6156 309454 -5536 344898
rect -6156 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 -5536 309454
rect -6156 309134 -5536 309218
rect -6156 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 -5536 309134
rect -6156 273454 -5536 308898
rect -6156 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 -5536 273454
rect -6156 273134 -5536 273218
rect -6156 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 -5536 273134
rect -6156 237454 -5536 272898
rect -6156 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 -5536 237454
rect -6156 237134 -5536 237218
rect -6156 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 -5536 237134
rect -6156 201454 -5536 236898
rect -6156 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 -5536 201454
rect -6156 201134 -5536 201218
rect -6156 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 -5536 201134
rect -6156 165454 -5536 200898
rect -6156 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 -5536 165454
rect -6156 165134 -5536 165218
rect -6156 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 -5536 165134
rect -6156 129454 -5536 164898
rect -6156 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 -5536 129454
rect -6156 129134 -5536 129218
rect -6156 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 -5536 129134
rect -6156 93454 -5536 128898
rect -6156 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 -5536 93454
rect -6156 93134 -5536 93218
rect -6156 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 -5536 93134
rect -6156 57454 -5536 92898
rect -6156 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 -5536 57454
rect -6156 57134 -5536 57218
rect -6156 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 -5536 57134
rect -6156 21454 -5536 56898
rect -6156 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 -5536 21454
rect -6156 21134 -5536 21218
rect -6156 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 -5536 21134
rect -6156 -4496 -5536 20898
rect -5196 708028 -4576 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 -4576 708028
rect -5196 707708 -4576 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 -4576 707708
rect -5196 700954 -4576 707472
rect -5196 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 -4576 700954
rect -5196 700634 -4576 700718
rect -5196 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 -4576 700634
rect -5196 664954 -4576 700398
rect -5196 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 -4576 664954
rect -5196 664634 -4576 664718
rect -5196 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 -4576 664634
rect -5196 628954 -4576 664398
rect -5196 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 -4576 628954
rect -5196 628634 -4576 628718
rect -5196 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 -4576 628634
rect -5196 592954 -4576 628398
rect -5196 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 -4576 592954
rect -5196 592634 -4576 592718
rect -5196 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 -4576 592634
rect -5196 556954 -4576 592398
rect -5196 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 -4576 556954
rect -5196 556634 -4576 556718
rect -5196 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 -4576 556634
rect -5196 520954 -4576 556398
rect -5196 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 -4576 520954
rect -5196 520634 -4576 520718
rect -5196 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 -4576 520634
rect -5196 484954 -4576 520398
rect -5196 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 -4576 484954
rect -5196 484634 -4576 484718
rect -5196 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 -4576 484634
rect -5196 448954 -4576 484398
rect -5196 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 -4576 448954
rect -5196 448634 -4576 448718
rect -5196 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 -4576 448634
rect -5196 412954 -4576 448398
rect -5196 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 -4576 412954
rect -5196 412634 -4576 412718
rect -5196 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 -4576 412634
rect -5196 376954 -4576 412398
rect -5196 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 -4576 376954
rect -5196 376634 -4576 376718
rect -5196 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 -4576 376634
rect -5196 340954 -4576 376398
rect -5196 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 -4576 340954
rect -5196 340634 -4576 340718
rect -5196 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 -4576 340634
rect -5196 304954 -4576 340398
rect -5196 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 -4576 304954
rect -5196 304634 -4576 304718
rect -5196 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 -4576 304634
rect -5196 268954 -4576 304398
rect -5196 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 -4576 268954
rect -5196 268634 -4576 268718
rect -5196 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 -4576 268634
rect -5196 232954 -4576 268398
rect -5196 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 -4576 232954
rect -5196 232634 -4576 232718
rect -5196 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 -4576 232634
rect -5196 196954 -4576 232398
rect -5196 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 -4576 196954
rect -5196 196634 -4576 196718
rect -5196 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 -4576 196634
rect -5196 160954 -4576 196398
rect -5196 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 -4576 160954
rect -5196 160634 -4576 160718
rect -5196 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 -4576 160634
rect -5196 124954 -4576 160398
rect -5196 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 -4576 124954
rect -5196 124634 -4576 124718
rect -5196 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 -4576 124634
rect -5196 88954 -4576 124398
rect -5196 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 -4576 88954
rect -5196 88634 -4576 88718
rect -5196 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 -4576 88634
rect -5196 52954 -4576 88398
rect -5196 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 -4576 52954
rect -5196 52634 -4576 52718
rect -5196 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 -4576 52634
rect -5196 16954 -4576 52398
rect -5196 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 -4576 16954
rect -5196 16634 -4576 16718
rect -5196 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 -4576 16634
rect -5196 -3536 -4576 16398
rect -4236 707068 -3616 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 -3616 707068
rect -4236 706748 -3616 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 -3616 706748
rect -4236 696454 -3616 706512
rect -4236 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 -3616 696454
rect -4236 696134 -3616 696218
rect -4236 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 -3616 696134
rect -4236 660454 -3616 695898
rect -4236 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 -3616 660454
rect -4236 660134 -3616 660218
rect -4236 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 -3616 660134
rect -4236 624454 -3616 659898
rect -4236 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 -3616 624454
rect -4236 624134 -3616 624218
rect -4236 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 -3616 624134
rect -4236 588454 -3616 623898
rect -4236 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 -3616 588454
rect -4236 588134 -3616 588218
rect -4236 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 -3616 588134
rect -4236 552454 -3616 587898
rect -4236 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 -3616 552454
rect -4236 552134 -3616 552218
rect -4236 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 -3616 552134
rect -4236 516454 -3616 551898
rect -4236 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 -3616 516454
rect -4236 516134 -3616 516218
rect -4236 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 -3616 516134
rect -4236 480454 -3616 515898
rect -4236 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 -3616 480454
rect -4236 480134 -3616 480218
rect -4236 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 -3616 480134
rect -4236 444454 -3616 479898
rect -4236 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 -3616 444454
rect -4236 444134 -3616 444218
rect -4236 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 -3616 444134
rect -4236 408454 -3616 443898
rect -4236 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 -3616 408454
rect -4236 408134 -3616 408218
rect -4236 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 -3616 408134
rect -4236 372454 -3616 407898
rect -4236 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 -3616 372454
rect -4236 372134 -3616 372218
rect -4236 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 -3616 372134
rect -4236 336454 -3616 371898
rect -4236 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 -3616 336454
rect -4236 336134 -3616 336218
rect -4236 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 -3616 336134
rect -4236 300454 -3616 335898
rect -4236 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 -3616 300454
rect -4236 300134 -3616 300218
rect -4236 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 -3616 300134
rect -4236 264454 -3616 299898
rect -4236 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 -3616 264454
rect -4236 264134 -3616 264218
rect -4236 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 -3616 264134
rect -4236 228454 -3616 263898
rect -4236 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 -3616 228454
rect -4236 228134 -3616 228218
rect -4236 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 -3616 228134
rect -4236 192454 -3616 227898
rect -4236 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 -3616 192454
rect -4236 192134 -3616 192218
rect -4236 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 -3616 192134
rect -4236 156454 -3616 191898
rect -4236 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 -3616 156454
rect -4236 156134 -3616 156218
rect -4236 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 -3616 156134
rect -4236 120454 -3616 155898
rect -4236 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 -3616 120454
rect -4236 120134 -3616 120218
rect -4236 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 -3616 120134
rect -4236 84454 -3616 119898
rect -4236 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 -3616 84454
rect -4236 84134 -3616 84218
rect -4236 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 -3616 84134
rect -4236 48454 -3616 83898
rect -4236 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 -3616 48454
rect -4236 48134 -3616 48218
rect -4236 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 -3616 48134
rect -4236 12454 -3616 47898
rect -4236 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 -3616 12454
rect -4236 12134 -3616 12218
rect -4236 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 -3616 12134
rect -4236 -2576 -3616 11898
rect -3276 706108 -2656 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 -2656 706108
rect -3276 705788 -2656 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 -2656 705788
rect -3276 691954 -2656 705552
rect -3276 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 -2656 691954
rect -3276 691634 -2656 691718
rect -3276 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 -2656 691634
rect -3276 655954 -2656 691398
rect -3276 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 -2656 655954
rect -3276 655634 -2656 655718
rect -3276 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 -2656 655634
rect -3276 619954 -2656 655398
rect -3276 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 -2656 619954
rect -3276 619634 -2656 619718
rect -3276 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 -2656 619634
rect -3276 583954 -2656 619398
rect -3276 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 -2656 583954
rect -3276 583634 -2656 583718
rect -3276 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 -2656 583634
rect -3276 547954 -2656 583398
rect -3276 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 -2656 547954
rect -3276 547634 -2656 547718
rect -3276 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 -2656 547634
rect -3276 511954 -2656 547398
rect -3276 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 -2656 511954
rect -3276 511634 -2656 511718
rect -3276 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 -2656 511634
rect -3276 475954 -2656 511398
rect -3276 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 -2656 475954
rect -3276 475634 -2656 475718
rect -3276 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 -2656 475634
rect -3276 439954 -2656 475398
rect -3276 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 -2656 439954
rect -3276 439634 -2656 439718
rect -3276 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 -2656 439634
rect -3276 403954 -2656 439398
rect -3276 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 -2656 403954
rect -3276 403634 -2656 403718
rect -3276 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 -2656 403634
rect -3276 367954 -2656 403398
rect -3276 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 -2656 367954
rect -3276 367634 -2656 367718
rect -3276 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 -2656 367634
rect -3276 331954 -2656 367398
rect -3276 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 -2656 331954
rect -3276 331634 -2656 331718
rect -3276 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 -2656 331634
rect -3276 295954 -2656 331398
rect -3276 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 -2656 295954
rect -3276 295634 -2656 295718
rect -3276 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 -2656 295634
rect -3276 259954 -2656 295398
rect -3276 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 -2656 259954
rect -3276 259634 -2656 259718
rect -3276 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 -2656 259634
rect -3276 223954 -2656 259398
rect -3276 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 -2656 223954
rect -3276 223634 -2656 223718
rect -3276 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 -2656 223634
rect -3276 187954 -2656 223398
rect -3276 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 -2656 187954
rect -3276 187634 -2656 187718
rect -3276 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 -2656 187634
rect -3276 151954 -2656 187398
rect -3276 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 -2656 151954
rect -3276 151634 -2656 151718
rect -3276 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 -2656 151634
rect -3276 115954 -2656 151398
rect -3276 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 -2656 115954
rect -3276 115634 -2656 115718
rect -3276 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 -2656 115634
rect -3276 79954 -2656 115398
rect -3276 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 -2656 79954
rect -3276 79634 -2656 79718
rect -3276 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 -2656 79634
rect -3276 43954 -2656 79398
rect -3276 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 -2656 43954
rect -3276 43634 -2656 43718
rect -3276 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 -2656 43634
rect -3276 7954 -2656 43398
rect -3276 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 -2656 7954
rect -3276 7634 -2656 7718
rect -3276 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 -2656 7634
rect -3276 -1616 -2656 7398
rect -2316 705148 -1696 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 -1696 705148
rect -2316 704828 -1696 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 -1696 704828
rect -2316 687454 -1696 704592
rect -2316 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 -1696 687454
rect -2316 687134 -1696 687218
rect -2316 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 -1696 687134
rect -2316 651454 -1696 686898
rect -2316 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 -1696 651454
rect -2316 651134 -1696 651218
rect -2316 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 -1696 651134
rect -2316 615454 -1696 650898
rect -2316 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 -1696 615454
rect -2316 615134 -1696 615218
rect -2316 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 -1696 615134
rect -2316 579454 -1696 614898
rect -2316 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 -1696 579454
rect -2316 579134 -1696 579218
rect -2316 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 -1696 579134
rect -2316 543454 -1696 578898
rect -2316 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 -1696 543454
rect -2316 543134 -1696 543218
rect -2316 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 -1696 543134
rect -2316 507454 -1696 542898
rect -2316 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 -1696 507454
rect -2316 507134 -1696 507218
rect -2316 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 -1696 507134
rect -2316 471454 -1696 506898
rect -2316 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 -1696 471454
rect -2316 471134 -1696 471218
rect -2316 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 -1696 471134
rect -2316 435454 -1696 470898
rect -2316 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 -1696 435454
rect -2316 435134 -1696 435218
rect -2316 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 -1696 435134
rect -2316 399454 -1696 434898
rect -2316 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 -1696 399454
rect -2316 399134 -1696 399218
rect -2316 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 -1696 399134
rect -2316 363454 -1696 398898
rect -2316 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 -1696 363454
rect -2316 363134 -1696 363218
rect -2316 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 -1696 363134
rect -2316 327454 -1696 362898
rect -2316 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 -1696 327454
rect -2316 327134 -1696 327218
rect -2316 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 -1696 327134
rect -2316 291454 -1696 326898
rect -2316 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 -1696 291454
rect -2316 291134 -1696 291218
rect -2316 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 -1696 291134
rect -2316 255454 -1696 290898
rect -2316 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 -1696 255454
rect -2316 255134 -1696 255218
rect -2316 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 -1696 255134
rect -2316 219454 -1696 254898
rect -2316 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 -1696 219454
rect -2316 219134 -1696 219218
rect -2316 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 -1696 219134
rect -2316 183454 -1696 218898
rect -2316 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 -1696 183454
rect -2316 183134 -1696 183218
rect -2316 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 -1696 183134
rect -2316 147454 -1696 182898
rect -2316 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 -1696 147454
rect -2316 147134 -1696 147218
rect -2316 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 -1696 147134
rect -2316 111454 -1696 146898
rect -2316 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 -1696 111454
rect -2316 111134 -1696 111218
rect -2316 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 -1696 111134
rect -2316 75454 -1696 110898
rect -2316 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 -1696 75454
rect -2316 75134 -1696 75218
rect -2316 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 -1696 75134
rect -2316 39454 -1696 74898
rect -2316 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 -1696 39454
rect -2316 39134 -1696 39218
rect -2316 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 -1696 39134
rect -2316 3454 -1696 38898
rect -2316 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 -1696 3454
rect -2316 3134 -1696 3218
rect -2316 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 -1696 3134
rect -2316 -656 -1696 2898
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 -1696 -656
rect -2316 -976 -1696 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 -1696 -976
rect -2316 -1244 -1696 -1212
rect 1794 705148 2414 711900
rect 1794 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 2414 705148
rect 1794 704828 2414 704912
rect 1794 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 2414 704828
rect 1794 687454 2414 704592
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -656 2414 2898
rect 1794 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 2414 -656
rect 1794 -976 2414 -892
rect 1794 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 2414 -976
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 -2656 -1616
rect -3276 -1936 -2656 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 -2656 -1936
rect -3276 -2204 -2656 -2172
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 -3616 -2576
rect -4236 -2896 -3616 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 -3616 -2896
rect -4236 -3164 -3616 -3132
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 -4576 -3536
rect -5196 -3856 -4576 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 -4576 -3856
rect -5196 -4124 -4576 -4092
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 -5536 -4496
rect -6156 -4816 -5536 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 -5536 -4816
rect -6156 -5084 -5536 -5052
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 -6496 -5456
rect -7116 -5776 -6496 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 -6496 -5776
rect -7116 -6044 -6496 -6012
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 -7456 -6416
rect -8076 -6736 -7456 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 -7456 -6736
rect -8076 -7004 -7456 -6972
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 -8416 -7376
rect -9036 -7696 -8416 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 -8416 -7696
rect -9036 -7964 -8416 -7932
rect 1794 -7964 2414 -1212
rect 6294 706108 6914 711900
rect 6294 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 6914 706108
rect 6294 705788 6914 705872
rect 6294 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 6914 705788
rect 6294 691954 6914 705552
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1616 6914 7398
rect 6294 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 6914 -1616
rect 6294 -1936 6914 -1852
rect 6294 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 6914 -1936
rect 6294 -7964 6914 -2172
rect 10794 707068 11414 711900
rect 10794 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 11414 707068
rect 10794 706748 11414 706832
rect 10794 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 11414 706748
rect 10794 696454 11414 706512
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2576 11414 11898
rect 10794 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 11414 -2576
rect 10794 -2896 11414 -2812
rect 10794 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 11414 -2896
rect 10794 -7964 11414 -3132
rect 15294 708028 15914 711900
rect 15294 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 15914 708028
rect 15294 707708 15914 707792
rect 15294 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 15914 707708
rect 15294 700954 15914 707472
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3536 15914 16398
rect 15294 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 15914 -3536
rect 15294 -3856 15914 -3772
rect 15294 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 15914 -3856
rect 15294 -7964 15914 -4092
rect 19794 708988 20414 711900
rect 19794 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 20414 708988
rect 19794 708668 20414 708752
rect 19794 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 20414 708668
rect 19794 669454 20414 708432
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4496 20414 20898
rect 19794 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 20414 -4496
rect 19794 -4816 20414 -4732
rect 19794 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 20414 -4816
rect 19794 -7964 20414 -5052
rect 24294 709948 24914 711900
rect 24294 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 24914 709948
rect 24294 709628 24914 709712
rect 24294 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 24914 709628
rect 24294 673954 24914 709392
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5456 24914 25398
rect 24294 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 24914 -5456
rect 24294 -5776 24914 -5692
rect 24294 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 24914 -5776
rect 24294 -7964 24914 -6012
rect 28794 710908 29414 711900
rect 28794 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 29414 710908
rect 28794 710588 29414 710672
rect 28794 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 29414 710588
rect 28794 678454 29414 710352
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6416 29414 29898
rect 28794 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 29414 -6416
rect 28794 -6736 29414 -6652
rect 28794 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 29414 -6736
rect 28794 -7964 29414 -6972
rect 33294 711868 33914 711900
rect 33294 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 33914 711868
rect 33294 711548 33914 711632
rect 33294 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 33914 711548
rect 33294 682954 33914 711312
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7376 33914 34398
rect 33294 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 33914 -7376
rect 33294 -7696 33914 -7612
rect 33294 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 33914 -7696
rect 33294 -7964 33914 -7932
rect 37794 705148 38414 711900
rect 37794 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 38414 705148
rect 37794 704828 38414 704912
rect 37794 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 38414 704828
rect 37794 687454 38414 704592
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -656 38414 2898
rect 37794 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 38414 -656
rect 37794 -976 38414 -892
rect 37794 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 38414 -976
rect 37794 -7964 38414 -1212
rect 42294 706108 42914 711900
rect 42294 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 42914 706108
rect 42294 705788 42914 705872
rect 42294 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 42914 705788
rect 42294 691954 42914 705552
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1616 42914 7398
rect 42294 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 42914 -1616
rect 42294 -1936 42914 -1852
rect 42294 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 42914 -1936
rect 42294 -7964 42914 -2172
rect 46794 707068 47414 711900
rect 46794 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 47414 707068
rect 46794 706748 47414 706832
rect 46794 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 47414 706748
rect 46794 696454 47414 706512
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2576 47414 11898
rect 46794 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 47414 -2576
rect 46794 -2896 47414 -2812
rect 46794 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 47414 -2896
rect 46794 -7964 47414 -3132
rect 51294 708028 51914 711900
rect 51294 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 51914 708028
rect 51294 707708 51914 707792
rect 51294 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 51914 707708
rect 51294 700954 51914 707472
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3536 51914 16398
rect 51294 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 51914 -3536
rect 51294 -3856 51914 -3772
rect 51294 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 51914 -3856
rect 51294 -7964 51914 -4092
rect 55794 708988 56414 711900
rect 55794 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 56414 708988
rect 55794 708668 56414 708752
rect 55794 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 56414 708668
rect 55794 669454 56414 708432
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4496 56414 20898
rect 55794 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 56414 -4496
rect 55794 -4816 56414 -4732
rect 55794 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 56414 -4816
rect 55794 -7964 56414 -5052
rect 60294 709948 60914 711900
rect 60294 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 60914 709948
rect 60294 709628 60914 709712
rect 60294 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 60914 709628
rect 60294 673954 60914 709392
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5456 60914 25398
rect 60294 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 60914 -5456
rect 60294 -5776 60914 -5692
rect 60294 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 60914 -5776
rect 60294 -7964 60914 -6012
rect 64794 710908 65414 711900
rect 64794 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 65414 710908
rect 64794 710588 65414 710672
rect 64794 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 65414 710588
rect 64794 678454 65414 710352
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6416 65414 29898
rect 64794 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 65414 -6416
rect 64794 -6736 65414 -6652
rect 64794 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 65414 -6736
rect 64794 -7964 65414 -6972
rect 69294 711868 69914 711900
rect 69294 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 69914 711868
rect 69294 711548 69914 711632
rect 69294 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 69914 711548
rect 69294 682954 69914 711312
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7376 69914 34398
rect 69294 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 69914 -7376
rect 69294 -7696 69914 -7612
rect 69294 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 69914 -7696
rect 69294 -7964 69914 -7932
rect 73794 705148 74414 711900
rect 73794 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 74414 705148
rect 73794 704828 74414 704912
rect 73794 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 74414 704828
rect 73794 687454 74414 704592
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -656 74414 2898
rect 73794 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 74414 -656
rect 73794 -976 74414 -892
rect 73794 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 74414 -976
rect 73794 -7964 74414 -1212
rect 78294 706108 78914 711900
rect 78294 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 78914 706108
rect 78294 705788 78914 705872
rect 78294 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 78914 705788
rect 78294 691954 78914 705552
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1616 78914 7398
rect 78294 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 78914 -1616
rect 78294 -1936 78914 -1852
rect 78294 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 78914 -1936
rect 78294 -7964 78914 -2172
rect 82794 707068 83414 711900
rect 82794 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 83414 707068
rect 82794 706748 83414 706832
rect 82794 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 83414 706748
rect 82794 696454 83414 706512
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2576 83414 11898
rect 82794 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 83414 -2576
rect 82794 -2896 83414 -2812
rect 82794 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 83414 -2896
rect 82794 -7964 83414 -3132
rect 87294 708028 87914 711900
rect 87294 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 87914 708028
rect 87294 707708 87914 707792
rect 87294 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 87914 707708
rect 87294 700954 87914 707472
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3536 87914 16398
rect 87294 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 87914 -3536
rect 87294 -3856 87914 -3772
rect 87294 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 87914 -3856
rect 87294 -7964 87914 -4092
rect 91794 708988 92414 711900
rect 91794 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 92414 708988
rect 91794 708668 92414 708752
rect 91794 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 92414 708668
rect 91794 669454 92414 708432
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4496 92414 20898
rect 91794 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 92414 -4496
rect 91794 -4816 92414 -4732
rect 91794 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 92414 -4816
rect 91794 -7964 92414 -5052
rect 96294 709948 96914 711900
rect 96294 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 96914 709948
rect 96294 709628 96914 709712
rect 96294 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 96914 709628
rect 96294 673954 96914 709392
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5456 96914 25398
rect 96294 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 96914 -5456
rect 96294 -5776 96914 -5692
rect 96294 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 96914 -5776
rect 96294 -7964 96914 -6012
rect 100794 710908 101414 711900
rect 100794 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 101414 710908
rect 100794 710588 101414 710672
rect 100794 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 101414 710588
rect 100794 678454 101414 710352
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6416 101414 29898
rect 100794 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 101414 -6416
rect 100794 -6736 101414 -6652
rect 100794 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 101414 -6736
rect 100794 -7964 101414 -6972
rect 105294 711868 105914 711900
rect 105294 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 105914 711868
rect 105294 711548 105914 711632
rect 105294 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 105914 711548
rect 105294 682954 105914 711312
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7376 105914 34398
rect 105294 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 105914 -7376
rect 105294 -7696 105914 -7612
rect 105294 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 105914 -7696
rect 105294 -7964 105914 -7932
rect 109794 705148 110414 711900
rect 109794 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 110414 705148
rect 109794 704828 110414 704912
rect 109794 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 110414 704828
rect 109794 687454 110414 704592
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -656 110414 2898
rect 109794 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 110414 -656
rect 109794 -976 110414 -892
rect 109794 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 110414 -976
rect 109794 -7964 110414 -1212
rect 114294 706108 114914 711900
rect 114294 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 114914 706108
rect 114294 705788 114914 705872
rect 114294 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 114914 705788
rect 114294 691954 114914 705552
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1616 114914 7398
rect 114294 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 114914 -1616
rect 114294 -1936 114914 -1852
rect 114294 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 114914 -1936
rect 114294 -7964 114914 -2172
rect 118794 707068 119414 711900
rect 118794 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 119414 707068
rect 118794 706748 119414 706832
rect 118794 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 119414 706748
rect 118794 696454 119414 706512
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2576 119414 11898
rect 118794 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 119414 -2576
rect 118794 -2896 119414 -2812
rect 118794 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 119414 -2896
rect 118794 -7964 119414 -3132
rect 123294 708028 123914 711900
rect 123294 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 123914 708028
rect 123294 707708 123914 707792
rect 123294 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 123914 707708
rect 123294 700954 123914 707472
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3536 123914 16398
rect 123294 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 123914 -3536
rect 123294 -3856 123914 -3772
rect 123294 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 123914 -3856
rect 123294 -7964 123914 -4092
rect 127794 708988 128414 711900
rect 127794 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 128414 708988
rect 127794 708668 128414 708752
rect 127794 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 128414 708668
rect 127794 669454 128414 708432
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4496 128414 20898
rect 127794 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 128414 -4496
rect 127794 -4816 128414 -4732
rect 127794 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 128414 -4816
rect 127794 -7964 128414 -5052
rect 132294 709948 132914 711900
rect 132294 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 132914 709948
rect 132294 709628 132914 709712
rect 132294 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 132914 709628
rect 132294 673954 132914 709392
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5456 132914 25398
rect 132294 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 132914 -5456
rect 132294 -5776 132914 -5692
rect 132294 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 132914 -5776
rect 132294 -7964 132914 -6012
rect 136794 710908 137414 711900
rect 136794 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 137414 710908
rect 136794 710588 137414 710672
rect 136794 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 137414 710588
rect 136794 678454 137414 710352
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6416 137414 29898
rect 136794 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 137414 -6416
rect 136794 -6736 137414 -6652
rect 136794 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 137414 -6736
rect 136794 -7964 137414 -6972
rect 141294 711868 141914 711900
rect 141294 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 141914 711868
rect 141294 711548 141914 711632
rect 141294 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 141914 711548
rect 141294 682954 141914 711312
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7376 141914 34398
rect 141294 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 141914 -7376
rect 141294 -7696 141914 -7612
rect 141294 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 141914 -7696
rect 141294 -7964 141914 -7932
rect 145794 705148 146414 711900
rect 145794 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 146414 705148
rect 145794 704828 146414 704912
rect 145794 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 146414 704828
rect 145794 687454 146414 704592
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -656 146414 2898
rect 145794 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 146414 -656
rect 145794 -976 146414 -892
rect 145794 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 146414 -976
rect 145794 -7964 146414 -1212
rect 150294 706108 150914 711900
rect 150294 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 150914 706108
rect 150294 705788 150914 705872
rect 150294 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 150914 705788
rect 150294 691954 150914 705552
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1616 150914 7398
rect 150294 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 150914 -1616
rect 150294 -1936 150914 -1852
rect 150294 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 150914 -1936
rect 150294 -7964 150914 -2172
rect 154794 707068 155414 711900
rect 154794 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 155414 707068
rect 154794 706748 155414 706832
rect 154794 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 155414 706748
rect 154794 696454 155414 706512
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2576 155414 11898
rect 154794 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 155414 -2576
rect 154794 -2896 155414 -2812
rect 154794 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 155414 -2896
rect 154794 -7964 155414 -3132
rect 159294 708028 159914 711900
rect 159294 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 159914 708028
rect 159294 707708 159914 707792
rect 159294 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 159914 707708
rect 159294 700954 159914 707472
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3536 159914 16398
rect 159294 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 159914 -3536
rect 159294 -3856 159914 -3772
rect 159294 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 159914 -3856
rect 159294 -7964 159914 -4092
rect 163794 708988 164414 711900
rect 163794 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 164414 708988
rect 163794 708668 164414 708752
rect 163794 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 164414 708668
rect 163794 669454 164414 708432
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4496 164414 20898
rect 163794 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 164414 -4496
rect 163794 -4816 164414 -4732
rect 163794 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 164414 -4816
rect 163794 -7964 164414 -5052
rect 168294 709948 168914 711900
rect 168294 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 168914 709948
rect 168294 709628 168914 709712
rect 168294 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 168914 709628
rect 168294 673954 168914 709392
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5456 168914 25398
rect 168294 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 168914 -5456
rect 168294 -5776 168914 -5692
rect 168294 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 168914 -5776
rect 168294 -7964 168914 -6012
rect 172794 710908 173414 711900
rect 172794 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 173414 710908
rect 172794 710588 173414 710672
rect 172794 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 173414 710588
rect 172794 678454 173414 710352
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6416 173414 29898
rect 172794 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 173414 -6416
rect 172794 -6736 173414 -6652
rect 172794 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 173414 -6736
rect 172794 -7964 173414 -6972
rect 177294 711868 177914 711900
rect 177294 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 177914 711868
rect 177294 711548 177914 711632
rect 177294 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 177914 711548
rect 177294 682954 177914 711312
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7376 177914 34398
rect 177294 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 177914 -7376
rect 177294 -7696 177914 -7612
rect 177294 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 177914 -7696
rect 177294 -7964 177914 -7932
rect 181794 705148 182414 711900
rect 181794 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 182414 705148
rect 181794 704828 182414 704912
rect 181794 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 182414 704828
rect 181794 687454 182414 704592
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -656 182414 2898
rect 181794 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 182414 -656
rect 181794 -976 182414 -892
rect 181794 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 182414 -976
rect 181794 -7964 182414 -1212
rect 186294 706108 186914 711900
rect 186294 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 186914 706108
rect 186294 705788 186914 705872
rect 186294 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 186914 705788
rect 186294 691954 186914 705552
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1616 186914 7398
rect 186294 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 186914 -1616
rect 186294 -1936 186914 -1852
rect 186294 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 186914 -1936
rect 186294 -7964 186914 -2172
rect 190794 707068 191414 711900
rect 190794 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 191414 707068
rect 190794 706748 191414 706832
rect 190794 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 191414 706748
rect 190794 696454 191414 706512
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2576 191414 11898
rect 190794 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 191414 -2576
rect 190794 -2896 191414 -2812
rect 190794 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 191414 -2896
rect 190794 -7964 191414 -3132
rect 195294 708028 195914 711900
rect 195294 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 195914 708028
rect 195294 707708 195914 707792
rect 195294 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 195914 707708
rect 195294 700954 195914 707472
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3536 195914 16398
rect 195294 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 195914 -3536
rect 195294 -3856 195914 -3772
rect 195294 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 195914 -3856
rect 195294 -7964 195914 -4092
rect 199794 708988 200414 711900
rect 199794 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 200414 708988
rect 199794 708668 200414 708752
rect 199794 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 200414 708668
rect 199794 669454 200414 708432
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4496 200414 20898
rect 199794 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 200414 -4496
rect 199794 -4816 200414 -4732
rect 199794 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 200414 -4816
rect 199794 -7964 200414 -5052
rect 204294 709948 204914 711900
rect 204294 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 204914 709948
rect 204294 709628 204914 709712
rect 204294 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 204914 709628
rect 204294 673954 204914 709392
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5456 204914 25398
rect 204294 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 204914 -5456
rect 204294 -5776 204914 -5692
rect 204294 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 204914 -5776
rect 204294 -7964 204914 -6012
rect 208794 710908 209414 711900
rect 208794 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 209414 710908
rect 208794 710588 209414 710672
rect 208794 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 209414 710588
rect 208794 678454 209414 710352
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6416 209414 29898
rect 208794 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 209414 -6416
rect 208794 -6736 209414 -6652
rect 208794 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 209414 -6736
rect 208794 -7964 209414 -6972
rect 213294 711868 213914 711900
rect 213294 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 213914 711868
rect 213294 711548 213914 711632
rect 213294 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 213914 711548
rect 213294 682954 213914 711312
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7376 213914 34398
rect 213294 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 213914 -7376
rect 213294 -7696 213914 -7612
rect 213294 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 213914 -7696
rect 213294 -7964 213914 -7932
rect 217794 705148 218414 711900
rect 217794 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 218414 705148
rect 217794 704828 218414 704912
rect 217794 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 218414 704828
rect 217794 687454 218414 704592
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -656 218414 2898
rect 217794 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 218414 -656
rect 217794 -976 218414 -892
rect 217794 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 218414 -976
rect 217794 -7964 218414 -1212
rect 222294 706108 222914 711900
rect 222294 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 222914 706108
rect 222294 705788 222914 705872
rect 222294 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 222914 705788
rect 222294 691954 222914 705552
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1616 222914 7398
rect 222294 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 222914 -1616
rect 222294 -1936 222914 -1852
rect 222294 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 222914 -1936
rect 222294 -7964 222914 -2172
rect 226794 707068 227414 711900
rect 226794 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 227414 707068
rect 226794 706748 227414 706832
rect 226794 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 227414 706748
rect 226794 696454 227414 706512
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 231294 708028 231914 711900
rect 231294 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 231914 708028
rect 231294 707708 231914 707792
rect 231294 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 231914 707708
rect 231294 700954 231914 707472
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 262000 231914 268398
rect 235794 708988 236414 711900
rect 235794 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 236414 708988
rect 235794 708668 236414 708752
rect 235794 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 236414 708668
rect 235794 669454 236414 708432
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 262000 236414 272898
rect 240294 709948 240914 711900
rect 240294 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 240914 709948
rect 240294 709628 240914 709712
rect 240294 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 240914 709628
rect 240294 673954 240914 709392
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 262000 240914 277398
rect 244794 710908 245414 711900
rect 244794 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 245414 710908
rect 244794 710588 245414 710672
rect 244794 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 245414 710588
rect 244794 678454 245414 710352
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 262000 245414 281898
rect 249294 711868 249914 711900
rect 249294 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 249914 711868
rect 249294 711548 249914 711632
rect 249294 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 249914 711548
rect 249294 682954 249914 711312
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 262000 249914 286398
rect 253794 705148 254414 711900
rect 253794 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 254414 705148
rect 253794 704828 254414 704912
rect 253794 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 254414 704828
rect 253794 687454 254414 704592
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 262000 254414 290898
rect 258294 706108 258914 711900
rect 258294 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 258914 706108
rect 258294 705788 258914 705872
rect 258294 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 258914 705788
rect 258294 691954 258914 705552
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 262000 258914 295398
rect 262794 707068 263414 711900
rect 262794 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 263414 707068
rect 262794 706748 263414 706832
rect 262794 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 263414 706748
rect 262794 696454 263414 706512
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 262000 263414 263898
rect 267294 708028 267914 711900
rect 267294 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 267914 708028
rect 267294 707708 267914 707792
rect 267294 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 267914 707708
rect 267294 700954 267914 707472
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 262000 267914 268398
rect 271794 708988 272414 711900
rect 271794 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 272414 708988
rect 271794 708668 272414 708752
rect 271794 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 272414 708668
rect 271794 669454 272414 708432
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 262000 272414 272898
rect 276294 709948 276914 711900
rect 276294 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 276914 709948
rect 276294 709628 276914 709712
rect 276294 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 276914 709628
rect 276294 673954 276914 709392
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 262000 276914 277398
rect 280794 710908 281414 711900
rect 280794 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 281414 710908
rect 280794 710588 281414 710672
rect 280794 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 281414 710588
rect 280794 678454 281414 710352
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 262000 281414 281898
rect 285294 711868 285914 711900
rect 285294 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 285914 711868
rect 285294 711548 285914 711632
rect 285294 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 285914 711548
rect 285294 682954 285914 711312
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 262000 285914 286398
rect 289794 705148 290414 711900
rect 289794 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 290414 705148
rect 289794 704828 290414 704912
rect 289794 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 290414 704828
rect 289794 687454 290414 704592
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 262000 290414 290898
rect 294294 706108 294914 711900
rect 294294 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 294914 706108
rect 294294 705788 294914 705872
rect 294294 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 294914 705788
rect 294294 691954 294914 705552
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 262000 294914 295398
rect 298794 707068 299414 711900
rect 298794 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 299414 707068
rect 298794 706748 299414 706832
rect 298794 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 299414 706748
rect 298794 696454 299414 706512
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 262000 299414 263898
rect 303294 708028 303914 711900
rect 303294 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 303914 708028
rect 303294 707708 303914 707792
rect 303294 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 303914 707708
rect 303294 700954 303914 707472
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 262000 303914 268398
rect 307794 708988 308414 711900
rect 307794 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 308414 708988
rect 307794 708668 308414 708752
rect 307794 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 308414 708668
rect 307794 669454 308414 708432
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 262000 308414 272898
rect 312294 709948 312914 711900
rect 312294 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 312914 709948
rect 312294 709628 312914 709712
rect 312294 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 312914 709628
rect 312294 673954 312914 709392
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 262000 312914 277398
rect 316794 710908 317414 711900
rect 316794 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 317414 710908
rect 316794 710588 317414 710672
rect 316794 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 317414 710588
rect 316794 678454 317414 710352
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 262000 317414 281898
rect 321294 711868 321914 711900
rect 321294 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 321914 711868
rect 321294 711548 321914 711632
rect 321294 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 321914 711548
rect 321294 682954 321914 711312
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 262000 321914 286398
rect 325794 705148 326414 711900
rect 325794 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 326414 705148
rect 325794 704828 326414 704912
rect 325794 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 326414 704828
rect 325794 687454 326414 704592
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 262000 326414 290898
rect 330294 706108 330914 711900
rect 330294 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 330914 706108
rect 330294 705788 330914 705872
rect 330294 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 330914 705788
rect 330294 691954 330914 705552
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 262000 330914 295398
rect 334794 707068 335414 711900
rect 334794 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 335414 707068
rect 334794 706748 335414 706832
rect 334794 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 335414 706748
rect 334794 696454 335414 706512
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 262000 335414 263898
rect 339294 708028 339914 711900
rect 339294 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 339914 708028
rect 339294 707708 339914 707792
rect 339294 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 339914 707708
rect 339294 700954 339914 707472
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 262000 339914 268398
rect 343794 708988 344414 711900
rect 343794 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 344414 708988
rect 343794 708668 344414 708752
rect 343794 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 344414 708668
rect 343794 669454 344414 708432
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 262000 344414 272898
rect 348294 709948 348914 711900
rect 348294 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 348914 709948
rect 348294 709628 348914 709712
rect 348294 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 348914 709628
rect 348294 673954 348914 709392
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 262000 348914 277398
rect 352794 710908 353414 711900
rect 352794 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 353414 710908
rect 352794 710588 353414 710672
rect 352794 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 353414 710588
rect 352794 678454 353414 710352
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 262000 353414 281898
rect 357294 711868 357914 711900
rect 357294 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 357914 711868
rect 357294 711548 357914 711632
rect 357294 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 357914 711548
rect 357294 682954 357914 711312
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 236208 255454 236528 255486
rect 236208 255218 236250 255454
rect 236486 255218 236528 255454
rect 236208 255134 236528 255218
rect 236208 254898 236250 255134
rect 236486 254898 236528 255134
rect 236208 254866 236528 254898
rect 266928 255454 267248 255486
rect 266928 255218 266970 255454
rect 267206 255218 267248 255454
rect 266928 255134 267248 255218
rect 266928 254898 266970 255134
rect 267206 254898 267248 255134
rect 266928 254866 267248 254898
rect 297648 255454 297968 255486
rect 297648 255218 297690 255454
rect 297926 255218 297968 255454
rect 297648 255134 297968 255218
rect 297648 254898 297690 255134
rect 297926 254898 297968 255134
rect 297648 254866 297968 254898
rect 328368 255454 328688 255486
rect 328368 255218 328410 255454
rect 328646 255218 328688 255454
rect 328368 255134 328688 255218
rect 328368 254898 328410 255134
rect 328646 254898 328688 255134
rect 328368 254866 328688 254898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 251568 223954 251888 223986
rect 251568 223718 251610 223954
rect 251846 223718 251888 223954
rect 251568 223634 251888 223718
rect 251568 223398 251610 223634
rect 251846 223398 251888 223634
rect 251568 223366 251888 223398
rect 282288 223954 282608 223986
rect 282288 223718 282330 223954
rect 282566 223718 282608 223954
rect 282288 223634 282608 223718
rect 282288 223398 282330 223634
rect 282566 223398 282608 223634
rect 282288 223366 282608 223398
rect 313008 223954 313328 223986
rect 313008 223718 313050 223954
rect 313286 223718 313328 223954
rect 313008 223634 313328 223718
rect 313008 223398 313050 223634
rect 313286 223398 313328 223634
rect 313008 223366 313328 223398
rect 343728 223954 344048 223986
rect 343728 223718 343770 223954
rect 344006 223718 344048 223954
rect 343728 223634 344048 223718
rect 343728 223398 343770 223634
rect 344006 223398 344048 223634
rect 343728 223366 344048 223398
rect 236208 219454 236528 219486
rect 236208 219218 236250 219454
rect 236486 219218 236528 219454
rect 236208 219134 236528 219218
rect 236208 218898 236250 219134
rect 236486 218898 236528 219134
rect 236208 218866 236528 218898
rect 266928 219454 267248 219486
rect 266928 219218 266970 219454
rect 267206 219218 267248 219454
rect 266928 219134 267248 219218
rect 266928 218898 266970 219134
rect 267206 218898 267248 219134
rect 266928 218866 267248 218898
rect 297648 219454 297968 219486
rect 297648 219218 297690 219454
rect 297926 219218 297968 219454
rect 297648 219134 297968 219218
rect 297648 218898 297690 219134
rect 297926 218898 297968 219134
rect 297648 218866 297968 218898
rect 328368 219454 328688 219486
rect 328368 219218 328410 219454
rect 328646 219218 328688 219454
rect 328368 219134 328688 219218
rect 328368 218898 328410 219134
rect 328646 218898 328688 219134
rect 328368 218866 328688 218898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 251568 187954 251888 187986
rect 251568 187718 251610 187954
rect 251846 187718 251888 187954
rect 251568 187634 251888 187718
rect 251568 187398 251610 187634
rect 251846 187398 251888 187634
rect 251568 187366 251888 187398
rect 282288 187954 282608 187986
rect 282288 187718 282330 187954
rect 282566 187718 282608 187954
rect 282288 187634 282608 187718
rect 282288 187398 282330 187634
rect 282566 187398 282608 187634
rect 282288 187366 282608 187398
rect 313008 187954 313328 187986
rect 313008 187718 313050 187954
rect 313286 187718 313328 187954
rect 313008 187634 313328 187718
rect 313008 187398 313050 187634
rect 313286 187398 313328 187634
rect 313008 187366 313328 187398
rect 343728 187954 344048 187986
rect 343728 187718 343770 187954
rect 344006 187718 344048 187954
rect 343728 187634 344048 187718
rect 343728 187398 343770 187634
rect 344006 187398 344048 187634
rect 343728 187366 344048 187398
rect 236208 183454 236528 183486
rect 236208 183218 236250 183454
rect 236486 183218 236528 183454
rect 236208 183134 236528 183218
rect 236208 182898 236250 183134
rect 236486 182898 236528 183134
rect 236208 182866 236528 182898
rect 266928 183454 267248 183486
rect 266928 183218 266970 183454
rect 267206 183218 267248 183454
rect 266928 183134 267248 183218
rect 266928 182898 266970 183134
rect 267206 182898 267248 183134
rect 266928 182866 267248 182898
rect 297648 183454 297968 183486
rect 297648 183218 297690 183454
rect 297926 183218 297968 183454
rect 297648 183134 297968 183218
rect 297648 182898 297690 183134
rect 297926 182898 297968 183134
rect 297648 182866 297968 182898
rect 328368 183454 328688 183486
rect 328368 183218 328410 183454
rect 328646 183218 328688 183454
rect 328368 183134 328688 183218
rect 328368 182898 328410 183134
rect 328646 182898 328688 183134
rect 328368 182866 328688 182898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 251568 151954 251888 151986
rect 251568 151718 251610 151954
rect 251846 151718 251888 151954
rect 251568 151634 251888 151718
rect 251568 151398 251610 151634
rect 251846 151398 251888 151634
rect 251568 151366 251888 151398
rect 282288 151954 282608 151986
rect 282288 151718 282330 151954
rect 282566 151718 282608 151954
rect 282288 151634 282608 151718
rect 282288 151398 282330 151634
rect 282566 151398 282608 151634
rect 282288 151366 282608 151398
rect 313008 151954 313328 151986
rect 313008 151718 313050 151954
rect 313286 151718 313328 151954
rect 313008 151634 313328 151718
rect 313008 151398 313050 151634
rect 313286 151398 313328 151634
rect 313008 151366 313328 151398
rect 343728 151954 344048 151986
rect 343728 151718 343770 151954
rect 344006 151718 344048 151954
rect 343728 151634 344048 151718
rect 343728 151398 343770 151634
rect 344006 151398 344048 151634
rect 343728 151366 344048 151398
rect 236208 147454 236528 147486
rect 236208 147218 236250 147454
rect 236486 147218 236528 147454
rect 236208 147134 236528 147218
rect 236208 146898 236250 147134
rect 236486 146898 236528 147134
rect 236208 146866 236528 146898
rect 266928 147454 267248 147486
rect 266928 147218 266970 147454
rect 267206 147218 267248 147454
rect 266928 147134 267248 147218
rect 266928 146898 266970 147134
rect 267206 146898 267248 147134
rect 266928 146866 267248 146898
rect 297648 147454 297968 147486
rect 297648 147218 297690 147454
rect 297926 147218 297968 147454
rect 297648 147134 297968 147218
rect 297648 146898 297690 147134
rect 297926 146898 297968 147134
rect 297648 146866 297968 146898
rect 328368 147454 328688 147486
rect 328368 147218 328410 147454
rect 328646 147218 328688 147454
rect 328368 147134 328688 147218
rect 328368 146898 328410 147134
rect 328646 146898 328688 147134
rect 328368 146866 328688 146898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 251568 115954 251888 115986
rect 251568 115718 251610 115954
rect 251846 115718 251888 115954
rect 251568 115634 251888 115718
rect 251568 115398 251610 115634
rect 251846 115398 251888 115634
rect 251568 115366 251888 115398
rect 282288 115954 282608 115986
rect 282288 115718 282330 115954
rect 282566 115718 282608 115954
rect 282288 115634 282608 115718
rect 282288 115398 282330 115634
rect 282566 115398 282608 115634
rect 282288 115366 282608 115398
rect 313008 115954 313328 115986
rect 313008 115718 313050 115954
rect 313286 115718 313328 115954
rect 313008 115634 313328 115718
rect 313008 115398 313050 115634
rect 313286 115398 313328 115634
rect 313008 115366 313328 115398
rect 343728 115954 344048 115986
rect 343728 115718 343770 115954
rect 344006 115718 344048 115954
rect 343728 115634 344048 115718
rect 343728 115398 343770 115634
rect 344006 115398 344048 115634
rect 343728 115366 344048 115398
rect 236208 111454 236528 111486
rect 236208 111218 236250 111454
rect 236486 111218 236528 111454
rect 236208 111134 236528 111218
rect 236208 110898 236250 111134
rect 236486 110898 236528 111134
rect 236208 110866 236528 110898
rect 266928 111454 267248 111486
rect 266928 111218 266970 111454
rect 267206 111218 267248 111454
rect 266928 111134 267248 111218
rect 266928 110898 266970 111134
rect 267206 110898 267248 111134
rect 266928 110866 267248 110898
rect 297648 111454 297968 111486
rect 297648 111218 297690 111454
rect 297926 111218 297968 111454
rect 297648 111134 297968 111218
rect 297648 110898 297690 111134
rect 297926 110898 297968 111134
rect 297648 110866 297968 110898
rect 328368 111454 328688 111486
rect 328368 111218 328410 111454
rect 328646 111218 328688 111454
rect 328368 111134 328688 111218
rect 328368 110898 328410 111134
rect 328646 110898 328688 111134
rect 328368 110866 328688 110898
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2576 227414 11898
rect 226794 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 227414 -2576
rect 226794 -2896 227414 -2812
rect 226794 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 227414 -2896
rect 226794 -7964 227414 -3132
rect 231294 88954 231914 98000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3536 231914 16398
rect 231294 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 231914 -3536
rect 231294 -3856 231914 -3772
rect 231294 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 231914 -3856
rect 231294 -7964 231914 -4092
rect 235794 93454 236414 98000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4496 236414 20898
rect 235794 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 236414 -4496
rect 235794 -4816 236414 -4732
rect 235794 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 236414 -4816
rect 235794 -7964 236414 -5052
rect 240294 97954 240914 98000
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5456 240914 25398
rect 240294 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 240914 -5456
rect 240294 -5776 240914 -5692
rect 240294 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 240914 -5776
rect 240294 -7964 240914 -6012
rect 244794 66454 245414 98000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6416 245414 29898
rect 244794 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 245414 -6416
rect 244794 -6736 245414 -6652
rect 244794 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 245414 -6736
rect 244794 -7964 245414 -6972
rect 249294 70954 249914 98000
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7376 249914 34398
rect 249294 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 249914 -7376
rect 249294 -7696 249914 -7612
rect 249294 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 249914 -7696
rect 249294 -7964 249914 -7932
rect 253794 75454 254414 98000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -656 254414 2898
rect 253794 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 254414 -656
rect 253794 -976 254414 -892
rect 253794 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 254414 -976
rect 253794 -7964 254414 -1212
rect 258294 79954 258914 98000
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1616 258914 7398
rect 258294 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 258914 -1616
rect 258294 -1936 258914 -1852
rect 258294 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 258914 -1936
rect 258294 -7964 258914 -2172
rect 262794 84454 263414 98000
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2576 263414 11898
rect 262794 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 263414 -2576
rect 262794 -2896 263414 -2812
rect 262794 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 263414 -2896
rect 262794 -7964 263414 -3132
rect 267294 88954 267914 98000
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3536 267914 16398
rect 267294 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 267914 -3536
rect 267294 -3856 267914 -3772
rect 267294 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 267914 -3856
rect 267294 -7964 267914 -4092
rect 271794 93454 272414 98000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4496 272414 20898
rect 271794 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 272414 -4496
rect 271794 -4816 272414 -4732
rect 271794 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 272414 -4816
rect 271794 -7964 272414 -5052
rect 276294 97954 276914 98000
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5456 276914 25398
rect 276294 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 276914 -5456
rect 276294 -5776 276914 -5692
rect 276294 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 276914 -5776
rect 276294 -7964 276914 -6012
rect 280794 66454 281414 98000
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6416 281414 29898
rect 280794 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 281414 -6416
rect 280794 -6736 281414 -6652
rect 280794 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 281414 -6736
rect 280794 -7964 281414 -6972
rect 285294 70954 285914 98000
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7376 285914 34398
rect 285294 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 285914 -7376
rect 285294 -7696 285914 -7612
rect 285294 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 285914 -7696
rect 285294 -7964 285914 -7932
rect 289794 75454 290414 98000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -656 290414 2898
rect 289794 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 290414 -656
rect 289794 -976 290414 -892
rect 289794 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 290414 -976
rect 289794 -7964 290414 -1212
rect 294294 79954 294914 98000
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1616 294914 7398
rect 294294 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 294914 -1616
rect 294294 -1936 294914 -1852
rect 294294 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 294914 -1936
rect 294294 -7964 294914 -2172
rect 298794 84454 299414 98000
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2576 299414 11898
rect 298794 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 299414 -2576
rect 298794 -2896 299414 -2812
rect 298794 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 299414 -2896
rect 298794 -7964 299414 -3132
rect 303294 88954 303914 98000
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3536 303914 16398
rect 303294 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 303914 -3536
rect 303294 -3856 303914 -3772
rect 303294 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 303914 -3856
rect 303294 -7964 303914 -4092
rect 307794 93454 308414 98000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4496 308414 20898
rect 307794 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 308414 -4496
rect 307794 -4816 308414 -4732
rect 307794 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 308414 -4816
rect 307794 -7964 308414 -5052
rect 312294 97954 312914 98000
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5456 312914 25398
rect 312294 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 312914 -5456
rect 312294 -5776 312914 -5692
rect 312294 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 312914 -5776
rect 312294 -7964 312914 -6012
rect 316794 66454 317414 98000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6416 317414 29898
rect 316794 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 317414 -6416
rect 316794 -6736 317414 -6652
rect 316794 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 317414 -6736
rect 316794 -7964 317414 -6972
rect 321294 70954 321914 98000
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7376 321914 34398
rect 321294 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 321914 -7376
rect 321294 -7696 321914 -7612
rect 321294 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 321914 -7696
rect 321294 -7964 321914 -7932
rect 325794 75454 326414 98000
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -656 326414 2898
rect 325794 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 326414 -656
rect 325794 -976 326414 -892
rect 325794 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 326414 -976
rect 325794 -7964 326414 -1212
rect 330294 79954 330914 98000
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1616 330914 7398
rect 330294 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 330914 -1616
rect 330294 -1936 330914 -1852
rect 330294 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 330914 -1936
rect 330294 -7964 330914 -2172
rect 334794 84454 335414 98000
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2576 335414 11898
rect 334794 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 335414 -2576
rect 334794 -2896 335414 -2812
rect 334794 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 335414 -2896
rect 334794 -7964 335414 -3132
rect 339294 88954 339914 98000
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3536 339914 16398
rect 339294 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 339914 -3536
rect 339294 -3856 339914 -3772
rect 339294 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 339914 -3856
rect 339294 -7964 339914 -4092
rect 343794 93454 344414 98000
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4496 344414 20898
rect 343794 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 344414 -4496
rect 343794 -4816 344414 -4732
rect 343794 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 344414 -4816
rect 343794 -7964 344414 -5052
rect 348294 97954 348914 98000
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5456 348914 25398
rect 348294 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 348914 -5456
rect 348294 -5776 348914 -5692
rect 348294 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 348914 -5776
rect 348294 -7964 348914 -6012
rect 352794 66454 353414 98000
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6416 353414 29898
rect 352794 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 353414 -6416
rect 352794 -6736 353414 -6652
rect 352794 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 353414 -6736
rect 352794 -7964 353414 -6972
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7376 357914 34398
rect 357294 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 357914 -7376
rect 357294 -7696 357914 -7612
rect 357294 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 357914 -7696
rect 357294 -7964 357914 -7932
rect 361794 705148 362414 711900
rect 361794 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 362414 705148
rect 361794 704828 362414 704912
rect 361794 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 362414 704828
rect 361794 687454 362414 704592
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -656 362414 2898
rect 361794 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 362414 -656
rect 361794 -976 362414 -892
rect 361794 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 362414 -976
rect 361794 -7964 362414 -1212
rect 366294 706108 366914 711900
rect 366294 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 366914 706108
rect 366294 705788 366914 705872
rect 366294 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 366914 705788
rect 366294 691954 366914 705552
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1616 366914 7398
rect 366294 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 366914 -1616
rect 366294 -1936 366914 -1852
rect 366294 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 366914 -1936
rect 366294 -7964 366914 -2172
rect 370794 707068 371414 711900
rect 370794 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 371414 707068
rect 370794 706748 371414 706832
rect 370794 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 371414 706748
rect 370794 696454 371414 706512
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2576 371414 11898
rect 370794 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 371414 -2576
rect 370794 -2896 371414 -2812
rect 370794 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 371414 -2896
rect 370794 -7964 371414 -3132
rect 375294 708028 375914 711900
rect 375294 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 375914 708028
rect 375294 707708 375914 707792
rect 375294 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 375914 707708
rect 375294 700954 375914 707472
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3536 375914 16398
rect 375294 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 375914 -3536
rect 375294 -3856 375914 -3772
rect 375294 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 375914 -3856
rect 375294 -7964 375914 -4092
rect 379794 708988 380414 711900
rect 379794 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 380414 708988
rect 379794 708668 380414 708752
rect 379794 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 380414 708668
rect 379794 669454 380414 708432
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4496 380414 20898
rect 379794 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 380414 -4496
rect 379794 -4816 380414 -4732
rect 379794 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 380414 -4816
rect 379794 -7964 380414 -5052
rect 384294 709948 384914 711900
rect 384294 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 384914 709948
rect 384294 709628 384914 709712
rect 384294 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 384914 709628
rect 384294 673954 384914 709392
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5456 384914 25398
rect 384294 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 384914 -5456
rect 384294 -5776 384914 -5692
rect 384294 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 384914 -5776
rect 384294 -7964 384914 -6012
rect 388794 710908 389414 711900
rect 388794 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 389414 710908
rect 388794 710588 389414 710672
rect 388794 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 389414 710588
rect 388794 678454 389414 710352
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6416 389414 29898
rect 388794 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 389414 -6416
rect 388794 -6736 389414 -6652
rect 388794 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 389414 -6736
rect 388794 -7964 389414 -6972
rect 393294 711868 393914 711900
rect 393294 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 393914 711868
rect 393294 711548 393914 711632
rect 393294 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 393914 711548
rect 393294 682954 393914 711312
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7376 393914 34398
rect 393294 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 393914 -7376
rect 393294 -7696 393914 -7612
rect 393294 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 393914 -7696
rect 393294 -7964 393914 -7932
rect 397794 705148 398414 711900
rect 397794 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 398414 705148
rect 397794 704828 398414 704912
rect 397794 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 398414 704828
rect 397794 687454 398414 704592
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -656 398414 2898
rect 397794 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 398414 -656
rect 397794 -976 398414 -892
rect 397794 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 398414 -976
rect 397794 -7964 398414 -1212
rect 402294 706108 402914 711900
rect 402294 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 402914 706108
rect 402294 705788 402914 705872
rect 402294 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 402914 705788
rect 402294 691954 402914 705552
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1616 402914 7398
rect 402294 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 402914 -1616
rect 402294 -1936 402914 -1852
rect 402294 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 402914 -1936
rect 402294 -7964 402914 -2172
rect 406794 707068 407414 711900
rect 406794 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 407414 707068
rect 406794 706748 407414 706832
rect 406794 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 407414 706748
rect 406794 696454 407414 706512
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2576 407414 11898
rect 406794 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 407414 -2576
rect 406794 -2896 407414 -2812
rect 406794 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 407414 -2896
rect 406794 -7964 407414 -3132
rect 411294 708028 411914 711900
rect 411294 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 411914 708028
rect 411294 707708 411914 707792
rect 411294 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 411914 707708
rect 411294 700954 411914 707472
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3536 411914 16398
rect 411294 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 411914 -3536
rect 411294 -3856 411914 -3772
rect 411294 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 411914 -3856
rect 411294 -7964 411914 -4092
rect 415794 708988 416414 711900
rect 415794 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 416414 708988
rect 415794 708668 416414 708752
rect 415794 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 416414 708668
rect 415794 669454 416414 708432
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4496 416414 20898
rect 415794 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 416414 -4496
rect 415794 -4816 416414 -4732
rect 415794 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 416414 -4816
rect 415794 -7964 416414 -5052
rect 420294 709948 420914 711900
rect 420294 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 420914 709948
rect 420294 709628 420914 709712
rect 420294 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 420914 709628
rect 420294 673954 420914 709392
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5456 420914 25398
rect 420294 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 420914 -5456
rect 420294 -5776 420914 -5692
rect 420294 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 420914 -5776
rect 420294 -7964 420914 -6012
rect 424794 710908 425414 711900
rect 424794 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 425414 710908
rect 424794 710588 425414 710672
rect 424794 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 425414 710588
rect 424794 678454 425414 710352
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6416 425414 29898
rect 424794 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 425414 -6416
rect 424794 -6736 425414 -6652
rect 424794 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 425414 -6736
rect 424794 -7964 425414 -6972
rect 429294 711868 429914 711900
rect 429294 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 429914 711868
rect 429294 711548 429914 711632
rect 429294 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 429914 711548
rect 429294 682954 429914 711312
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7376 429914 34398
rect 429294 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 429914 -7376
rect 429294 -7696 429914 -7612
rect 429294 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 429914 -7696
rect 429294 -7964 429914 -7932
rect 433794 705148 434414 711900
rect 433794 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 434414 705148
rect 433794 704828 434414 704912
rect 433794 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 434414 704828
rect 433794 687454 434414 704592
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -656 434414 2898
rect 433794 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 434414 -656
rect 433794 -976 434414 -892
rect 433794 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 434414 -976
rect 433794 -7964 434414 -1212
rect 438294 706108 438914 711900
rect 438294 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 438914 706108
rect 438294 705788 438914 705872
rect 438294 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 438914 705788
rect 438294 691954 438914 705552
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1616 438914 7398
rect 438294 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 438914 -1616
rect 438294 -1936 438914 -1852
rect 438294 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 438914 -1936
rect 438294 -7964 438914 -2172
rect 442794 707068 443414 711900
rect 442794 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 443414 707068
rect 442794 706748 443414 706832
rect 442794 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 443414 706748
rect 442794 696454 443414 706512
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2576 443414 11898
rect 442794 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 443414 -2576
rect 442794 -2896 443414 -2812
rect 442794 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 443414 -2896
rect 442794 -7964 443414 -3132
rect 447294 708028 447914 711900
rect 447294 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 447914 708028
rect 447294 707708 447914 707792
rect 447294 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 447914 707708
rect 447294 700954 447914 707472
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3536 447914 16398
rect 447294 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 447914 -3536
rect 447294 -3856 447914 -3772
rect 447294 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 447914 -3856
rect 447294 -7964 447914 -4092
rect 451794 708988 452414 711900
rect 451794 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 452414 708988
rect 451794 708668 452414 708752
rect 451794 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 452414 708668
rect 451794 669454 452414 708432
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4496 452414 20898
rect 451794 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 452414 -4496
rect 451794 -4816 452414 -4732
rect 451794 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 452414 -4816
rect 451794 -7964 452414 -5052
rect 456294 709948 456914 711900
rect 456294 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 456914 709948
rect 456294 709628 456914 709712
rect 456294 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 456914 709628
rect 456294 673954 456914 709392
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5456 456914 25398
rect 456294 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 456914 -5456
rect 456294 -5776 456914 -5692
rect 456294 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 456914 -5776
rect 456294 -7964 456914 -6012
rect 460794 710908 461414 711900
rect 460794 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 461414 710908
rect 460794 710588 461414 710672
rect 460794 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 461414 710588
rect 460794 678454 461414 710352
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6416 461414 29898
rect 460794 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 461414 -6416
rect 460794 -6736 461414 -6652
rect 460794 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 461414 -6736
rect 460794 -7964 461414 -6972
rect 465294 711868 465914 711900
rect 465294 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 465914 711868
rect 465294 711548 465914 711632
rect 465294 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 465914 711548
rect 465294 682954 465914 711312
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7376 465914 34398
rect 465294 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 465914 -7376
rect 465294 -7696 465914 -7612
rect 465294 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 465914 -7696
rect 465294 -7964 465914 -7932
rect 469794 705148 470414 711900
rect 469794 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 470414 705148
rect 469794 704828 470414 704912
rect 469794 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 470414 704828
rect 469794 687454 470414 704592
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -656 470414 2898
rect 469794 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 470414 -656
rect 469794 -976 470414 -892
rect 469794 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 470414 -976
rect 469794 -7964 470414 -1212
rect 474294 706108 474914 711900
rect 474294 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 474914 706108
rect 474294 705788 474914 705872
rect 474294 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 474914 705788
rect 474294 691954 474914 705552
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1616 474914 7398
rect 474294 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 474914 -1616
rect 474294 -1936 474914 -1852
rect 474294 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 474914 -1936
rect 474294 -7964 474914 -2172
rect 478794 707068 479414 711900
rect 478794 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 479414 707068
rect 478794 706748 479414 706832
rect 478794 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 479414 706748
rect 478794 696454 479414 706512
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2576 479414 11898
rect 478794 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 479414 -2576
rect 478794 -2896 479414 -2812
rect 478794 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 479414 -2896
rect 478794 -7964 479414 -3132
rect 483294 708028 483914 711900
rect 483294 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 483914 708028
rect 483294 707708 483914 707792
rect 483294 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 483914 707708
rect 483294 700954 483914 707472
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3536 483914 16398
rect 483294 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 483914 -3536
rect 483294 -3856 483914 -3772
rect 483294 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 483914 -3856
rect 483294 -7964 483914 -4092
rect 487794 708988 488414 711900
rect 487794 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 488414 708988
rect 487794 708668 488414 708752
rect 487794 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 488414 708668
rect 487794 669454 488414 708432
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4496 488414 20898
rect 487794 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 488414 -4496
rect 487794 -4816 488414 -4732
rect 487794 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 488414 -4816
rect 487794 -7964 488414 -5052
rect 492294 709948 492914 711900
rect 492294 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 492914 709948
rect 492294 709628 492914 709712
rect 492294 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 492914 709628
rect 492294 673954 492914 709392
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5456 492914 25398
rect 492294 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 492914 -5456
rect 492294 -5776 492914 -5692
rect 492294 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 492914 -5776
rect 492294 -7964 492914 -6012
rect 496794 710908 497414 711900
rect 496794 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 497414 710908
rect 496794 710588 497414 710672
rect 496794 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 497414 710588
rect 496794 678454 497414 710352
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6416 497414 29898
rect 496794 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 497414 -6416
rect 496794 -6736 497414 -6652
rect 496794 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 497414 -6736
rect 496794 -7964 497414 -6972
rect 501294 711868 501914 711900
rect 501294 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 501914 711868
rect 501294 711548 501914 711632
rect 501294 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 501914 711548
rect 501294 682954 501914 711312
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7376 501914 34398
rect 501294 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 501914 -7376
rect 501294 -7696 501914 -7612
rect 501294 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 501914 -7696
rect 501294 -7964 501914 -7932
rect 505794 705148 506414 711900
rect 505794 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 506414 705148
rect 505794 704828 506414 704912
rect 505794 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 506414 704828
rect 505794 687454 506414 704592
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -656 506414 2898
rect 505794 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 506414 -656
rect 505794 -976 506414 -892
rect 505794 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 506414 -976
rect 505794 -7964 506414 -1212
rect 510294 706108 510914 711900
rect 510294 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 510914 706108
rect 510294 705788 510914 705872
rect 510294 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 510914 705788
rect 510294 691954 510914 705552
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1616 510914 7398
rect 510294 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 510914 -1616
rect 510294 -1936 510914 -1852
rect 510294 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 510914 -1936
rect 510294 -7964 510914 -2172
rect 514794 707068 515414 711900
rect 514794 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 515414 707068
rect 514794 706748 515414 706832
rect 514794 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 515414 706748
rect 514794 696454 515414 706512
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2576 515414 11898
rect 514794 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 515414 -2576
rect 514794 -2896 515414 -2812
rect 514794 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 515414 -2896
rect 514794 -7964 515414 -3132
rect 519294 708028 519914 711900
rect 519294 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 519914 708028
rect 519294 707708 519914 707792
rect 519294 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 519914 707708
rect 519294 700954 519914 707472
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3536 519914 16398
rect 519294 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 519914 -3536
rect 519294 -3856 519914 -3772
rect 519294 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 519914 -3856
rect 519294 -7964 519914 -4092
rect 523794 708988 524414 711900
rect 523794 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 524414 708988
rect 523794 708668 524414 708752
rect 523794 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 524414 708668
rect 523794 669454 524414 708432
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4496 524414 20898
rect 523794 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 524414 -4496
rect 523794 -4816 524414 -4732
rect 523794 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 524414 -4816
rect 523794 -7964 524414 -5052
rect 528294 709948 528914 711900
rect 528294 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 528914 709948
rect 528294 709628 528914 709712
rect 528294 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 528914 709628
rect 528294 673954 528914 709392
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5456 528914 25398
rect 528294 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 528914 -5456
rect 528294 -5776 528914 -5692
rect 528294 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 528914 -5776
rect 528294 -7964 528914 -6012
rect 532794 710908 533414 711900
rect 532794 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 533414 710908
rect 532794 710588 533414 710672
rect 532794 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 533414 710588
rect 532794 678454 533414 710352
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6416 533414 29898
rect 532794 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 533414 -6416
rect 532794 -6736 533414 -6652
rect 532794 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 533414 -6736
rect 532794 -7964 533414 -6972
rect 537294 711868 537914 711900
rect 537294 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 537914 711868
rect 537294 711548 537914 711632
rect 537294 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 537914 711548
rect 537294 682954 537914 711312
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7376 537914 34398
rect 537294 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 537914 -7376
rect 537294 -7696 537914 -7612
rect 537294 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 537914 -7696
rect 537294 -7964 537914 -7932
rect 541794 705148 542414 711900
rect 541794 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 542414 705148
rect 541794 704828 542414 704912
rect 541794 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 542414 704828
rect 541794 687454 542414 704592
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -656 542414 2898
rect 541794 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 542414 -656
rect 541794 -976 542414 -892
rect 541794 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 542414 -976
rect 541794 -7964 542414 -1212
rect 546294 706108 546914 711900
rect 546294 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 546914 706108
rect 546294 705788 546914 705872
rect 546294 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 546914 705788
rect 546294 691954 546914 705552
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1616 546914 7398
rect 546294 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 546914 -1616
rect 546294 -1936 546914 -1852
rect 546294 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 546914 -1936
rect 546294 -7964 546914 -2172
rect 550794 707068 551414 711900
rect 550794 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 551414 707068
rect 550794 706748 551414 706832
rect 550794 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 551414 706748
rect 550794 696454 551414 706512
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2576 551414 11898
rect 550794 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 551414 -2576
rect 550794 -2896 551414 -2812
rect 550794 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 551414 -2896
rect 550794 -7964 551414 -3132
rect 555294 708028 555914 711900
rect 555294 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 555914 708028
rect 555294 707708 555914 707792
rect 555294 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 555914 707708
rect 555294 700954 555914 707472
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3536 555914 16398
rect 555294 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 555914 -3536
rect 555294 -3856 555914 -3772
rect 555294 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 555914 -3856
rect 555294 -7964 555914 -4092
rect 559794 708988 560414 711900
rect 559794 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 560414 708988
rect 559794 708668 560414 708752
rect 559794 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 560414 708668
rect 559794 669454 560414 708432
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4496 560414 20898
rect 559794 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 560414 -4496
rect 559794 -4816 560414 -4732
rect 559794 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 560414 -4816
rect 559794 -7964 560414 -5052
rect 564294 709948 564914 711900
rect 564294 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 564914 709948
rect 564294 709628 564914 709712
rect 564294 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 564914 709628
rect 564294 673954 564914 709392
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5456 564914 25398
rect 564294 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 564914 -5456
rect 564294 -5776 564914 -5692
rect 564294 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 564914 -5776
rect 564294 -7964 564914 -6012
rect 568794 710908 569414 711900
rect 568794 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 569414 710908
rect 568794 710588 569414 710672
rect 568794 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 569414 710588
rect 568794 678454 569414 710352
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6416 569414 29898
rect 568794 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 569414 -6416
rect 568794 -6736 569414 -6652
rect 568794 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 569414 -6736
rect 568794 -7964 569414 -6972
rect 573294 711868 573914 711900
rect 573294 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 573914 711868
rect 573294 711548 573914 711632
rect 573294 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 573914 711548
rect 573294 682954 573914 711312
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7376 573914 34398
rect 573294 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 573914 -7376
rect 573294 -7696 573914 -7612
rect 573294 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 573914 -7696
rect 573294 -7964 573914 -7932
rect 577794 705148 578414 711900
rect 577794 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 578414 705148
rect 577794 704828 578414 704912
rect 577794 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 578414 704828
rect 577794 687454 578414 704592
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -656 578414 2898
rect 577794 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 578414 -656
rect 577794 -976 578414 -892
rect 577794 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 578414 -976
rect 577794 -7964 578414 -1212
rect 582294 706108 582914 711900
rect 592340 711868 592960 711900
rect 592340 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect 592340 711548 592960 711632
rect 592340 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect 591380 710908 592000 710940
rect 591380 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect 591380 710588 592000 710672
rect 591380 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect 590420 709948 591040 709980
rect 590420 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect 590420 709628 591040 709712
rect 590420 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect 589460 708988 590080 709020
rect 589460 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect 589460 708668 590080 708752
rect 589460 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect 588500 708028 589120 708060
rect 588500 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect 588500 707708 589120 707792
rect 588500 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect 587540 707068 588160 707100
rect 587540 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect 587540 706748 588160 706832
rect 587540 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect 582294 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 582914 706108
rect 582294 705788 582914 705872
rect 582294 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 582914 705788
rect 582294 691954 582914 705552
rect 586580 706108 587200 706140
rect 586580 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect 586580 705788 587200 705872
rect 586580 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1616 582914 7398
rect 585620 705148 586240 705180
rect 585620 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect 585620 704828 586240 704912
rect 585620 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect 585620 687454 586240 704592
rect 585620 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 586240 687454
rect 585620 687134 586240 687218
rect 585620 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 586240 687134
rect 585620 651454 586240 686898
rect 585620 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 586240 651454
rect 585620 651134 586240 651218
rect 585620 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 586240 651134
rect 585620 615454 586240 650898
rect 585620 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 586240 615454
rect 585620 615134 586240 615218
rect 585620 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 586240 615134
rect 585620 579454 586240 614898
rect 585620 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 586240 579454
rect 585620 579134 586240 579218
rect 585620 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 586240 579134
rect 585620 543454 586240 578898
rect 585620 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 586240 543454
rect 585620 543134 586240 543218
rect 585620 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 586240 543134
rect 585620 507454 586240 542898
rect 585620 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 586240 507454
rect 585620 507134 586240 507218
rect 585620 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 586240 507134
rect 585620 471454 586240 506898
rect 585620 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 586240 471454
rect 585620 471134 586240 471218
rect 585620 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 586240 471134
rect 585620 435454 586240 470898
rect 585620 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 586240 435454
rect 585620 435134 586240 435218
rect 585620 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 586240 435134
rect 585620 399454 586240 434898
rect 585620 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 586240 399454
rect 585620 399134 586240 399218
rect 585620 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 586240 399134
rect 585620 363454 586240 398898
rect 585620 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 586240 363454
rect 585620 363134 586240 363218
rect 585620 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 586240 363134
rect 585620 327454 586240 362898
rect 585620 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 586240 327454
rect 585620 327134 586240 327218
rect 585620 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 586240 327134
rect 585620 291454 586240 326898
rect 585620 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 586240 291454
rect 585620 291134 586240 291218
rect 585620 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 586240 291134
rect 585620 255454 586240 290898
rect 585620 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 586240 255454
rect 585620 255134 586240 255218
rect 585620 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 586240 255134
rect 585620 219454 586240 254898
rect 585620 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 586240 219454
rect 585620 219134 586240 219218
rect 585620 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 586240 219134
rect 585620 183454 586240 218898
rect 585620 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 586240 183454
rect 585620 183134 586240 183218
rect 585620 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 586240 183134
rect 585620 147454 586240 182898
rect 585620 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 586240 147454
rect 585620 147134 586240 147218
rect 585620 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 586240 147134
rect 585620 111454 586240 146898
rect 585620 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 586240 111454
rect 585620 111134 586240 111218
rect 585620 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 586240 111134
rect 585620 75454 586240 110898
rect 585620 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 586240 75454
rect 585620 75134 586240 75218
rect 585620 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 586240 75134
rect 585620 39454 586240 74898
rect 585620 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 586240 39454
rect 585620 39134 586240 39218
rect 585620 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 586240 39134
rect 585620 3454 586240 38898
rect 585620 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 586240 3454
rect 585620 3134 586240 3218
rect 585620 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 586240 3134
rect 585620 -656 586240 2898
rect 585620 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect 585620 -976 586240 -892
rect 585620 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect 585620 -1244 586240 -1212
rect 586580 691954 587200 705552
rect 586580 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 587200 691954
rect 586580 691634 587200 691718
rect 586580 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 587200 691634
rect 586580 655954 587200 691398
rect 586580 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 587200 655954
rect 586580 655634 587200 655718
rect 586580 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 587200 655634
rect 586580 619954 587200 655398
rect 586580 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 587200 619954
rect 586580 619634 587200 619718
rect 586580 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 587200 619634
rect 586580 583954 587200 619398
rect 586580 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 587200 583954
rect 586580 583634 587200 583718
rect 586580 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 587200 583634
rect 586580 547954 587200 583398
rect 586580 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 587200 547954
rect 586580 547634 587200 547718
rect 586580 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 587200 547634
rect 586580 511954 587200 547398
rect 586580 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 587200 511954
rect 586580 511634 587200 511718
rect 586580 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 587200 511634
rect 586580 475954 587200 511398
rect 586580 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 587200 475954
rect 586580 475634 587200 475718
rect 586580 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 587200 475634
rect 586580 439954 587200 475398
rect 586580 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 587200 439954
rect 586580 439634 587200 439718
rect 586580 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 587200 439634
rect 586580 403954 587200 439398
rect 586580 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 587200 403954
rect 586580 403634 587200 403718
rect 586580 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 587200 403634
rect 586580 367954 587200 403398
rect 586580 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 587200 367954
rect 586580 367634 587200 367718
rect 586580 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 587200 367634
rect 586580 331954 587200 367398
rect 586580 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 587200 331954
rect 586580 331634 587200 331718
rect 586580 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 587200 331634
rect 586580 295954 587200 331398
rect 586580 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 587200 295954
rect 586580 295634 587200 295718
rect 586580 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 587200 295634
rect 586580 259954 587200 295398
rect 586580 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 587200 259954
rect 586580 259634 587200 259718
rect 586580 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 587200 259634
rect 586580 223954 587200 259398
rect 586580 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 587200 223954
rect 586580 223634 587200 223718
rect 586580 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 587200 223634
rect 586580 187954 587200 223398
rect 586580 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 587200 187954
rect 586580 187634 587200 187718
rect 586580 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 587200 187634
rect 586580 151954 587200 187398
rect 586580 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 587200 151954
rect 586580 151634 587200 151718
rect 586580 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 587200 151634
rect 586580 115954 587200 151398
rect 586580 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 587200 115954
rect 586580 115634 587200 115718
rect 586580 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 587200 115634
rect 586580 79954 587200 115398
rect 586580 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 587200 79954
rect 586580 79634 587200 79718
rect 586580 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 587200 79634
rect 586580 43954 587200 79398
rect 586580 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 587200 43954
rect 586580 43634 587200 43718
rect 586580 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 587200 43634
rect 586580 7954 587200 43398
rect 586580 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 587200 7954
rect 586580 7634 587200 7718
rect 586580 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 587200 7634
rect 582294 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 582914 -1616
rect 582294 -1936 582914 -1852
rect 582294 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 582914 -1936
rect 582294 -7964 582914 -2172
rect 586580 -1616 587200 7398
rect 586580 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect 586580 -1936 587200 -1852
rect 586580 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect 586580 -2204 587200 -2172
rect 587540 696454 588160 706512
rect 587540 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 588160 696454
rect 587540 696134 588160 696218
rect 587540 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 588160 696134
rect 587540 660454 588160 695898
rect 587540 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 588160 660454
rect 587540 660134 588160 660218
rect 587540 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 588160 660134
rect 587540 624454 588160 659898
rect 587540 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 588160 624454
rect 587540 624134 588160 624218
rect 587540 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 588160 624134
rect 587540 588454 588160 623898
rect 587540 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 588160 588454
rect 587540 588134 588160 588218
rect 587540 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 588160 588134
rect 587540 552454 588160 587898
rect 587540 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 588160 552454
rect 587540 552134 588160 552218
rect 587540 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 588160 552134
rect 587540 516454 588160 551898
rect 587540 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 588160 516454
rect 587540 516134 588160 516218
rect 587540 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 588160 516134
rect 587540 480454 588160 515898
rect 587540 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 588160 480454
rect 587540 480134 588160 480218
rect 587540 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 588160 480134
rect 587540 444454 588160 479898
rect 587540 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 588160 444454
rect 587540 444134 588160 444218
rect 587540 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 588160 444134
rect 587540 408454 588160 443898
rect 587540 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 588160 408454
rect 587540 408134 588160 408218
rect 587540 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 588160 408134
rect 587540 372454 588160 407898
rect 587540 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 588160 372454
rect 587540 372134 588160 372218
rect 587540 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 588160 372134
rect 587540 336454 588160 371898
rect 587540 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 588160 336454
rect 587540 336134 588160 336218
rect 587540 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 588160 336134
rect 587540 300454 588160 335898
rect 587540 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 588160 300454
rect 587540 300134 588160 300218
rect 587540 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 588160 300134
rect 587540 264454 588160 299898
rect 587540 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 588160 264454
rect 587540 264134 588160 264218
rect 587540 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 588160 264134
rect 587540 228454 588160 263898
rect 587540 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 588160 228454
rect 587540 228134 588160 228218
rect 587540 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 588160 228134
rect 587540 192454 588160 227898
rect 587540 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 588160 192454
rect 587540 192134 588160 192218
rect 587540 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 588160 192134
rect 587540 156454 588160 191898
rect 587540 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 588160 156454
rect 587540 156134 588160 156218
rect 587540 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 588160 156134
rect 587540 120454 588160 155898
rect 587540 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 588160 120454
rect 587540 120134 588160 120218
rect 587540 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 588160 120134
rect 587540 84454 588160 119898
rect 587540 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 588160 84454
rect 587540 84134 588160 84218
rect 587540 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 588160 84134
rect 587540 48454 588160 83898
rect 587540 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 588160 48454
rect 587540 48134 588160 48218
rect 587540 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 588160 48134
rect 587540 12454 588160 47898
rect 587540 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 588160 12454
rect 587540 12134 588160 12218
rect 587540 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 588160 12134
rect 587540 -2576 588160 11898
rect 587540 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect 587540 -2896 588160 -2812
rect 587540 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect 587540 -3164 588160 -3132
rect 588500 700954 589120 707472
rect 588500 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 589120 700954
rect 588500 700634 589120 700718
rect 588500 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 589120 700634
rect 588500 664954 589120 700398
rect 588500 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 589120 664954
rect 588500 664634 589120 664718
rect 588500 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 589120 664634
rect 588500 628954 589120 664398
rect 588500 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 589120 628954
rect 588500 628634 589120 628718
rect 588500 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 589120 628634
rect 588500 592954 589120 628398
rect 588500 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 589120 592954
rect 588500 592634 589120 592718
rect 588500 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 589120 592634
rect 588500 556954 589120 592398
rect 588500 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 589120 556954
rect 588500 556634 589120 556718
rect 588500 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 589120 556634
rect 588500 520954 589120 556398
rect 588500 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 589120 520954
rect 588500 520634 589120 520718
rect 588500 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 589120 520634
rect 588500 484954 589120 520398
rect 588500 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 589120 484954
rect 588500 484634 589120 484718
rect 588500 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 589120 484634
rect 588500 448954 589120 484398
rect 588500 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 589120 448954
rect 588500 448634 589120 448718
rect 588500 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 589120 448634
rect 588500 412954 589120 448398
rect 588500 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 589120 412954
rect 588500 412634 589120 412718
rect 588500 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 589120 412634
rect 588500 376954 589120 412398
rect 588500 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 589120 376954
rect 588500 376634 589120 376718
rect 588500 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 589120 376634
rect 588500 340954 589120 376398
rect 588500 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 589120 340954
rect 588500 340634 589120 340718
rect 588500 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 589120 340634
rect 588500 304954 589120 340398
rect 588500 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 589120 304954
rect 588500 304634 589120 304718
rect 588500 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 589120 304634
rect 588500 268954 589120 304398
rect 588500 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 589120 268954
rect 588500 268634 589120 268718
rect 588500 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 589120 268634
rect 588500 232954 589120 268398
rect 588500 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 589120 232954
rect 588500 232634 589120 232718
rect 588500 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 589120 232634
rect 588500 196954 589120 232398
rect 588500 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 589120 196954
rect 588500 196634 589120 196718
rect 588500 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 589120 196634
rect 588500 160954 589120 196398
rect 588500 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 589120 160954
rect 588500 160634 589120 160718
rect 588500 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 589120 160634
rect 588500 124954 589120 160398
rect 588500 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 589120 124954
rect 588500 124634 589120 124718
rect 588500 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 589120 124634
rect 588500 88954 589120 124398
rect 588500 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 589120 88954
rect 588500 88634 589120 88718
rect 588500 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 589120 88634
rect 588500 52954 589120 88398
rect 588500 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 589120 52954
rect 588500 52634 589120 52718
rect 588500 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 589120 52634
rect 588500 16954 589120 52398
rect 588500 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 589120 16954
rect 588500 16634 589120 16718
rect 588500 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 589120 16634
rect 588500 -3536 589120 16398
rect 588500 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect 588500 -3856 589120 -3772
rect 588500 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect 588500 -4124 589120 -4092
rect 589460 669454 590080 708432
rect 589460 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 590080 669454
rect 589460 669134 590080 669218
rect 589460 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 590080 669134
rect 589460 633454 590080 668898
rect 589460 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 590080 633454
rect 589460 633134 590080 633218
rect 589460 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 590080 633134
rect 589460 597454 590080 632898
rect 589460 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 590080 597454
rect 589460 597134 590080 597218
rect 589460 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 590080 597134
rect 589460 561454 590080 596898
rect 589460 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 590080 561454
rect 589460 561134 590080 561218
rect 589460 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 590080 561134
rect 589460 525454 590080 560898
rect 589460 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 590080 525454
rect 589460 525134 590080 525218
rect 589460 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 590080 525134
rect 589460 489454 590080 524898
rect 589460 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 590080 489454
rect 589460 489134 590080 489218
rect 589460 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 590080 489134
rect 589460 453454 590080 488898
rect 589460 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 590080 453454
rect 589460 453134 590080 453218
rect 589460 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 590080 453134
rect 589460 417454 590080 452898
rect 589460 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 590080 417454
rect 589460 417134 590080 417218
rect 589460 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 590080 417134
rect 589460 381454 590080 416898
rect 589460 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 590080 381454
rect 589460 381134 590080 381218
rect 589460 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 590080 381134
rect 589460 345454 590080 380898
rect 589460 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 590080 345454
rect 589460 345134 590080 345218
rect 589460 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 590080 345134
rect 589460 309454 590080 344898
rect 589460 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 590080 309454
rect 589460 309134 590080 309218
rect 589460 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 590080 309134
rect 589460 273454 590080 308898
rect 589460 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 590080 273454
rect 589460 273134 590080 273218
rect 589460 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 590080 273134
rect 589460 237454 590080 272898
rect 589460 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 590080 237454
rect 589460 237134 590080 237218
rect 589460 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 590080 237134
rect 589460 201454 590080 236898
rect 589460 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 590080 201454
rect 589460 201134 590080 201218
rect 589460 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 590080 201134
rect 589460 165454 590080 200898
rect 589460 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 590080 165454
rect 589460 165134 590080 165218
rect 589460 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 590080 165134
rect 589460 129454 590080 164898
rect 589460 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 590080 129454
rect 589460 129134 590080 129218
rect 589460 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 590080 129134
rect 589460 93454 590080 128898
rect 589460 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 590080 93454
rect 589460 93134 590080 93218
rect 589460 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 590080 93134
rect 589460 57454 590080 92898
rect 589460 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 590080 57454
rect 589460 57134 590080 57218
rect 589460 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 590080 57134
rect 589460 21454 590080 56898
rect 589460 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 590080 21454
rect 589460 21134 590080 21218
rect 589460 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 590080 21134
rect 589460 -4496 590080 20898
rect 589460 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect 589460 -4816 590080 -4732
rect 589460 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect 589460 -5084 590080 -5052
rect 590420 673954 591040 709392
rect 590420 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 591040 673954
rect 590420 673634 591040 673718
rect 590420 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 591040 673634
rect 590420 637954 591040 673398
rect 590420 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 591040 637954
rect 590420 637634 591040 637718
rect 590420 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 591040 637634
rect 590420 601954 591040 637398
rect 590420 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 591040 601954
rect 590420 601634 591040 601718
rect 590420 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 591040 601634
rect 590420 565954 591040 601398
rect 590420 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 591040 565954
rect 590420 565634 591040 565718
rect 590420 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 591040 565634
rect 590420 529954 591040 565398
rect 590420 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 591040 529954
rect 590420 529634 591040 529718
rect 590420 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 591040 529634
rect 590420 493954 591040 529398
rect 590420 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 591040 493954
rect 590420 493634 591040 493718
rect 590420 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 591040 493634
rect 590420 457954 591040 493398
rect 590420 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 591040 457954
rect 590420 457634 591040 457718
rect 590420 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 591040 457634
rect 590420 421954 591040 457398
rect 590420 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 591040 421954
rect 590420 421634 591040 421718
rect 590420 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 591040 421634
rect 590420 385954 591040 421398
rect 590420 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 591040 385954
rect 590420 385634 591040 385718
rect 590420 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 591040 385634
rect 590420 349954 591040 385398
rect 590420 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 591040 349954
rect 590420 349634 591040 349718
rect 590420 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 591040 349634
rect 590420 313954 591040 349398
rect 590420 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 591040 313954
rect 590420 313634 591040 313718
rect 590420 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 591040 313634
rect 590420 277954 591040 313398
rect 590420 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 591040 277954
rect 590420 277634 591040 277718
rect 590420 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 591040 277634
rect 590420 241954 591040 277398
rect 590420 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 591040 241954
rect 590420 241634 591040 241718
rect 590420 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 591040 241634
rect 590420 205954 591040 241398
rect 590420 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 591040 205954
rect 590420 205634 591040 205718
rect 590420 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 591040 205634
rect 590420 169954 591040 205398
rect 590420 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 591040 169954
rect 590420 169634 591040 169718
rect 590420 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 591040 169634
rect 590420 133954 591040 169398
rect 590420 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 591040 133954
rect 590420 133634 591040 133718
rect 590420 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 591040 133634
rect 590420 97954 591040 133398
rect 590420 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 591040 97954
rect 590420 97634 591040 97718
rect 590420 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 591040 97634
rect 590420 61954 591040 97398
rect 590420 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 591040 61954
rect 590420 61634 591040 61718
rect 590420 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 591040 61634
rect 590420 25954 591040 61398
rect 590420 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 591040 25954
rect 590420 25634 591040 25718
rect 590420 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 591040 25634
rect 590420 -5456 591040 25398
rect 590420 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect 590420 -5776 591040 -5692
rect 590420 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect 590420 -6044 591040 -6012
rect 591380 678454 592000 710352
rect 591380 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592000 678454
rect 591380 678134 592000 678218
rect 591380 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592000 678134
rect 591380 642454 592000 677898
rect 591380 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592000 642454
rect 591380 642134 592000 642218
rect 591380 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592000 642134
rect 591380 606454 592000 641898
rect 591380 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592000 606454
rect 591380 606134 592000 606218
rect 591380 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592000 606134
rect 591380 570454 592000 605898
rect 591380 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592000 570454
rect 591380 570134 592000 570218
rect 591380 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592000 570134
rect 591380 534454 592000 569898
rect 591380 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592000 534454
rect 591380 534134 592000 534218
rect 591380 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592000 534134
rect 591380 498454 592000 533898
rect 591380 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592000 498454
rect 591380 498134 592000 498218
rect 591380 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592000 498134
rect 591380 462454 592000 497898
rect 591380 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592000 462454
rect 591380 462134 592000 462218
rect 591380 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592000 462134
rect 591380 426454 592000 461898
rect 591380 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592000 426454
rect 591380 426134 592000 426218
rect 591380 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592000 426134
rect 591380 390454 592000 425898
rect 591380 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592000 390454
rect 591380 390134 592000 390218
rect 591380 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592000 390134
rect 591380 354454 592000 389898
rect 591380 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592000 354454
rect 591380 354134 592000 354218
rect 591380 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592000 354134
rect 591380 318454 592000 353898
rect 591380 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592000 318454
rect 591380 318134 592000 318218
rect 591380 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592000 318134
rect 591380 282454 592000 317898
rect 591380 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592000 282454
rect 591380 282134 592000 282218
rect 591380 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592000 282134
rect 591380 246454 592000 281898
rect 591380 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592000 246454
rect 591380 246134 592000 246218
rect 591380 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592000 246134
rect 591380 210454 592000 245898
rect 591380 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592000 210454
rect 591380 210134 592000 210218
rect 591380 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592000 210134
rect 591380 174454 592000 209898
rect 591380 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592000 174454
rect 591380 174134 592000 174218
rect 591380 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592000 174134
rect 591380 138454 592000 173898
rect 591380 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592000 138454
rect 591380 138134 592000 138218
rect 591380 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592000 138134
rect 591380 102454 592000 137898
rect 591380 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592000 102454
rect 591380 102134 592000 102218
rect 591380 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592000 102134
rect 591380 66454 592000 101898
rect 591380 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592000 66454
rect 591380 66134 592000 66218
rect 591380 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592000 66134
rect 591380 30454 592000 65898
rect 591380 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592000 30454
rect 591380 30134 592000 30218
rect 591380 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592000 30134
rect 591380 -6416 592000 29898
rect 591380 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect 591380 -6736 592000 -6652
rect 591380 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect 591380 -7004 592000 -6972
rect 592340 682954 592960 711312
rect 592340 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect 592340 682634 592960 682718
rect 592340 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect 592340 646954 592960 682398
rect 592340 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect 592340 646634 592960 646718
rect 592340 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect 592340 610954 592960 646398
rect 592340 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect 592340 610634 592960 610718
rect 592340 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect 592340 574954 592960 610398
rect 592340 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect 592340 574634 592960 574718
rect 592340 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect 592340 538954 592960 574398
rect 592340 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect 592340 538634 592960 538718
rect 592340 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect 592340 502954 592960 538398
rect 592340 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect 592340 502634 592960 502718
rect 592340 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect 592340 466954 592960 502398
rect 592340 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect 592340 466634 592960 466718
rect 592340 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect 592340 430954 592960 466398
rect 592340 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect 592340 430634 592960 430718
rect 592340 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect 592340 394954 592960 430398
rect 592340 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect 592340 394634 592960 394718
rect 592340 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect 592340 358954 592960 394398
rect 592340 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect 592340 358634 592960 358718
rect 592340 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect 592340 322954 592960 358398
rect 592340 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect 592340 322634 592960 322718
rect 592340 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect 592340 286954 592960 322398
rect 592340 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect 592340 286634 592960 286718
rect 592340 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect 592340 250954 592960 286398
rect 592340 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect 592340 250634 592960 250718
rect 592340 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect 592340 214954 592960 250398
rect 592340 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect 592340 214634 592960 214718
rect 592340 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect 592340 178954 592960 214398
rect 592340 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect 592340 178634 592960 178718
rect 592340 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect 592340 142954 592960 178398
rect 592340 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect 592340 142634 592960 142718
rect 592340 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect 592340 106954 592960 142398
rect 592340 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect 592340 106634 592960 106718
rect 592340 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect 592340 70954 592960 106398
rect 592340 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect 592340 70634 592960 70718
rect 592340 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect 592340 34954 592960 70398
rect 592340 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect 592340 34634 592960 34718
rect 592340 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect 592340 -7376 592960 34398
rect 592340 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect 592340 -7696 592960 -7612
rect 592340 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect 592340 -7964 592960 -7932
<< via4 >>
rect -9004 711632 -8768 711868
rect -8684 711632 -8448 711868
rect -9004 711312 -8768 711548
rect -8684 711312 -8448 711548
rect -9004 682718 -8768 682954
rect -8684 682718 -8448 682954
rect -9004 682398 -8768 682634
rect -8684 682398 -8448 682634
rect -9004 646718 -8768 646954
rect -8684 646718 -8448 646954
rect -9004 646398 -8768 646634
rect -8684 646398 -8448 646634
rect -9004 610718 -8768 610954
rect -8684 610718 -8448 610954
rect -9004 610398 -8768 610634
rect -8684 610398 -8448 610634
rect -9004 574718 -8768 574954
rect -8684 574718 -8448 574954
rect -9004 574398 -8768 574634
rect -8684 574398 -8448 574634
rect -9004 538718 -8768 538954
rect -8684 538718 -8448 538954
rect -9004 538398 -8768 538634
rect -8684 538398 -8448 538634
rect -9004 502718 -8768 502954
rect -8684 502718 -8448 502954
rect -9004 502398 -8768 502634
rect -8684 502398 -8448 502634
rect -9004 466718 -8768 466954
rect -8684 466718 -8448 466954
rect -9004 466398 -8768 466634
rect -8684 466398 -8448 466634
rect -9004 430718 -8768 430954
rect -8684 430718 -8448 430954
rect -9004 430398 -8768 430634
rect -8684 430398 -8448 430634
rect -9004 394718 -8768 394954
rect -8684 394718 -8448 394954
rect -9004 394398 -8768 394634
rect -8684 394398 -8448 394634
rect -9004 358718 -8768 358954
rect -8684 358718 -8448 358954
rect -9004 358398 -8768 358634
rect -8684 358398 -8448 358634
rect -9004 322718 -8768 322954
rect -8684 322718 -8448 322954
rect -9004 322398 -8768 322634
rect -8684 322398 -8448 322634
rect -9004 286718 -8768 286954
rect -8684 286718 -8448 286954
rect -9004 286398 -8768 286634
rect -8684 286398 -8448 286634
rect -9004 250718 -8768 250954
rect -8684 250718 -8448 250954
rect -9004 250398 -8768 250634
rect -8684 250398 -8448 250634
rect -9004 214718 -8768 214954
rect -8684 214718 -8448 214954
rect -9004 214398 -8768 214634
rect -8684 214398 -8448 214634
rect -9004 178718 -8768 178954
rect -8684 178718 -8448 178954
rect -9004 178398 -8768 178634
rect -8684 178398 -8448 178634
rect -9004 142718 -8768 142954
rect -8684 142718 -8448 142954
rect -9004 142398 -8768 142634
rect -8684 142398 -8448 142634
rect -9004 106718 -8768 106954
rect -8684 106718 -8448 106954
rect -9004 106398 -8768 106634
rect -8684 106398 -8448 106634
rect -9004 70718 -8768 70954
rect -8684 70718 -8448 70954
rect -9004 70398 -8768 70634
rect -8684 70398 -8448 70634
rect -9004 34718 -8768 34954
rect -8684 34718 -8448 34954
rect -9004 34398 -8768 34634
rect -8684 34398 -8448 34634
rect -8044 710672 -7808 710908
rect -7724 710672 -7488 710908
rect -8044 710352 -7808 710588
rect -7724 710352 -7488 710588
rect -8044 678218 -7808 678454
rect -7724 678218 -7488 678454
rect -8044 677898 -7808 678134
rect -7724 677898 -7488 678134
rect -8044 642218 -7808 642454
rect -7724 642218 -7488 642454
rect -8044 641898 -7808 642134
rect -7724 641898 -7488 642134
rect -8044 606218 -7808 606454
rect -7724 606218 -7488 606454
rect -8044 605898 -7808 606134
rect -7724 605898 -7488 606134
rect -8044 570218 -7808 570454
rect -7724 570218 -7488 570454
rect -8044 569898 -7808 570134
rect -7724 569898 -7488 570134
rect -8044 534218 -7808 534454
rect -7724 534218 -7488 534454
rect -8044 533898 -7808 534134
rect -7724 533898 -7488 534134
rect -8044 498218 -7808 498454
rect -7724 498218 -7488 498454
rect -8044 497898 -7808 498134
rect -7724 497898 -7488 498134
rect -8044 462218 -7808 462454
rect -7724 462218 -7488 462454
rect -8044 461898 -7808 462134
rect -7724 461898 -7488 462134
rect -8044 426218 -7808 426454
rect -7724 426218 -7488 426454
rect -8044 425898 -7808 426134
rect -7724 425898 -7488 426134
rect -8044 390218 -7808 390454
rect -7724 390218 -7488 390454
rect -8044 389898 -7808 390134
rect -7724 389898 -7488 390134
rect -8044 354218 -7808 354454
rect -7724 354218 -7488 354454
rect -8044 353898 -7808 354134
rect -7724 353898 -7488 354134
rect -8044 318218 -7808 318454
rect -7724 318218 -7488 318454
rect -8044 317898 -7808 318134
rect -7724 317898 -7488 318134
rect -8044 282218 -7808 282454
rect -7724 282218 -7488 282454
rect -8044 281898 -7808 282134
rect -7724 281898 -7488 282134
rect -8044 246218 -7808 246454
rect -7724 246218 -7488 246454
rect -8044 245898 -7808 246134
rect -7724 245898 -7488 246134
rect -8044 210218 -7808 210454
rect -7724 210218 -7488 210454
rect -8044 209898 -7808 210134
rect -7724 209898 -7488 210134
rect -8044 174218 -7808 174454
rect -7724 174218 -7488 174454
rect -8044 173898 -7808 174134
rect -7724 173898 -7488 174134
rect -8044 138218 -7808 138454
rect -7724 138218 -7488 138454
rect -8044 137898 -7808 138134
rect -7724 137898 -7488 138134
rect -8044 102218 -7808 102454
rect -7724 102218 -7488 102454
rect -8044 101898 -7808 102134
rect -7724 101898 -7488 102134
rect -8044 66218 -7808 66454
rect -7724 66218 -7488 66454
rect -8044 65898 -7808 66134
rect -7724 65898 -7488 66134
rect -8044 30218 -7808 30454
rect -7724 30218 -7488 30454
rect -8044 29898 -7808 30134
rect -7724 29898 -7488 30134
rect -7084 709712 -6848 709948
rect -6764 709712 -6528 709948
rect -7084 709392 -6848 709628
rect -6764 709392 -6528 709628
rect -7084 673718 -6848 673954
rect -6764 673718 -6528 673954
rect -7084 673398 -6848 673634
rect -6764 673398 -6528 673634
rect -7084 637718 -6848 637954
rect -6764 637718 -6528 637954
rect -7084 637398 -6848 637634
rect -6764 637398 -6528 637634
rect -7084 601718 -6848 601954
rect -6764 601718 -6528 601954
rect -7084 601398 -6848 601634
rect -6764 601398 -6528 601634
rect -7084 565718 -6848 565954
rect -6764 565718 -6528 565954
rect -7084 565398 -6848 565634
rect -6764 565398 -6528 565634
rect -7084 529718 -6848 529954
rect -6764 529718 -6528 529954
rect -7084 529398 -6848 529634
rect -6764 529398 -6528 529634
rect -7084 493718 -6848 493954
rect -6764 493718 -6528 493954
rect -7084 493398 -6848 493634
rect -6764 493398 -6528 493634
rect -7084 457718 -6848 457954
rect -6764 457718 -6528 457954
rect -7084 457398 -6848 457634
rect -6764 457398 -6528 457634
rect -7084 421718 -6848 421954
rect -6764 421718 -6528 421954
rect -7084 421398 -6848 421634
rect -6764 421398 -6528 421634
rect -7084 385718 -6848 385954
rect -6764 385718 -6528 385954
rect -7084 385398 -6848 385634
rect -6764 385398 -6528 385634
rect -7084 349718 -6848 349954
rect -6764 349718 -6528 349954
rect -7084 349398 -6848 349634
rect -6764 349398 -6528 349634
rect -7084 313718 -6848 313954
rect -6764 313718 -6528 313954
rect -7084 313398 -6848 313634
rect -6764 313398 -6528 313634
rect -7084 277718 -6848 277954
rect -6764 277718 -6528 277954
rect -7084 277398 -6848 277634
rect -6764 277398 -6528 277634
rect -7084 241718 -6848 241954
rect -6764 241718 -6528 241954
rect -7084 241398 -6848 241634
rect -6764 241398 -6528 241634
rect -7084 205718 -6848 205954
rect -6764 205718 -6528 205954
rect -7084 205398 -6848 205634
rect -6764 205398 -6528 205634
rect -7084 169718 -6848 169954
rect -6764 169718 -6528 169954
rect -7084 169398 -6848 169634
rect -6764 169398 -6528 169634
rect -7084 133718 -6848 133954
rect -6764 133718 -6528 133954
rect -7084 133398 -6848 133634
rect -6764 133398 -6528 133634
rect -7084 97718 -6848 97954
rect -6764 97718 -6528 97954
rect -7084 97398 -6848 97634
rect -6764 97398 -6528 97634
rect -7084 61718 -6848 61954
rect -6764 61718 -6528 61954
rect -7084 61398 -6848 61634
rect -6764 61398 -6528 61634
rect -7084 25718 -6848 25954
rect -6764 25718 -6528 25954
rect -7084 25398 -6848 25634
rect -6764 25398 -6528 25634
rect -6124 708752 -5888 708988
rect -5804 708752 -5568 708988
rect -6124 708432 -5888 708668
rect -5804 708432 -5568 708668
rect -6124 669218 -5888 669454
rect -5804 669218 -5568 669454
rect -6124 668898 -5888 669134
rect -5804 668898 -5568 669134
rect -6124 633218 -5888 633454
rect -5804 633218 -5568 633454
rect -6124 632898 -5888 633134
rect -5804 632898 -5568 633134
rect -6124 597218 -5888 597454
rect -5804 597218 -5568 597454
rect -6124 596898 -5888 597134
rect -5804 596898 -5568 597134
rect -6124 561218 -5888 561454
rect -5804 561218 -5568 561454
rect -6124 560898 -5888 561134
rect -5804 560898 -5568 561134
rect -6124 525218 -5888 525454
rect -5804 525218 -5568 525454
rect -6124 524898 -5888 525134
rect -5804 524898 -5568 525134
rect -6124 489218 -5888 489454
rect -5804 489218 -5568 489454
rect -6124 488898 -5888 489134
rect -5804 488898 -5568 489134
rect -6124 453218 -5888 453454
rect -5804 453218 -5568 453454
rect -6124 452898 -5888 453134
rect -5804 452898 -5568 453134
rect -6124 417218 -5888 417454
rect -5804 417218 -5568 417454
rect -6124 416898 -5888 417134
rect -5804 416898 -5568 417134
rect -6124 381218 -5888 381454
rect -5804 381218 -5568 381454
rect -6124 380898 -5888 381134
rect -5804 380898 -5568 381134
rect -6124 345218 -5888 345454
rect -5804 345218 -5568 345454
rect -6124 344898 -5888 345134
rect -5804 344898 -5568 345134
rect -6124 309218 -5888 309454
rect -5804 309218 -5568 309454
rect -6124 308898 -5888 309134
rect -5804 308898 -5568 309134
rect -6124 273218 -5888 273454
rect -5804 273218 -5568 273454
rect -6124 272898 -5888 273134
rect -5804 272898 -5568 273134
rect -6124 237218 -5888 237454
rect -5804 237218 -5568 237454
rect -6124 236898 -5888 237134
rect -5804 236898 -5568 237134
rect -6124 201218 -5888 201454
rect -5804 201218 -5568 201454
rect -6124 200898 -5888 201134
rect -5804 200898 -5568 201134
rect -6124 165218 -5888 165454
rect -5804 165218 -5568 165454
rect -6124 164898 -5888 165134
rect -5804 164898 -5568 165134
rect -6124 129218 -5888 129454
rect -5804 129218 -5568 129454
rect -6124 128898 -5888 129134
rect -5804 128898 -5568 129134
rect -6124 93218 -5888 93454
rect -5804 93218 -5568 93454
rect -6124 92898 -5888 93134
rect -5804 92898 -5568 93134
rect -6124 57218 -5888 57454
rect -5804 57218 -5568 57454
rect -6124 56898 -5888 57134
rect -5804 56898 -5568 57134
rect -6124 21218 -5888 21454
rect -5804 21218 -5568 21454
rect -6124 20898 -5888 21134
rect -5804 20898 -5568 21134
rect -5164 707792 -4928 708028
rect -4844 707792 -4608 708028
rect -5164 707472 -4928 707708
rect -4844 707472 -4608 707708
rect -5164 700718 -4928 700954
rect -4844 700718 -4608 700954
rect -5164 700398 -4928 700634
rect -4844 700398 -4608 700634
rect -5164 664718 -4928 664954
rect -4844 664718 -4608 664954
rect -5164 664398 -4928 664634
rect -4844 664398 -4608 664634
rect -5164 628718 -4928 628954
rect -4844 628718 -4608 628954
rect -5164 628398 -4928 628634
rect -4844 628398 -4608 628634
rect -5164 592718 -4928 592954
rect -4844 592718 -4608 592954
rect -5164 592398 -4928 592634
rect -4844 592398 -4608 592634
rect -5164 556718 -4928 556954
rect -4844 556718 -4608 556954
rect -5164 556398 -4928 556634
rect -4844 556398 -4608 556634
rect -5164 520718 -4928 520954
rect -4844 520718 -4608 520954
rect -5164 520398 -4928 520634
rect -4844 520398 -4608 520634
rect -5164 484718 -4928 484954
rect -4844 484718 -4608 484954
rect -5164 484398 -4928 484634
rect -4844 484398 -4608 484634
rect -5164 448718 -4928 448954
rect -4844 448718 -4608 448954
rect -5164 448398 -4928 448634
rect -4844 448398 -4608 448634
rect -5164 412718 -4928 412954
rect -4844 412718 -4608 412954
rect -5164 412398 -4928 412634
rect -4844 412398 -4608 412634
rect -5164 376718 -4928 376954
rect -4844 376718 -4608 376954
rect -5164 376398 -4928 376634
rect -4844 376398 -4608 376634
rect -5164 340718 -4928 340954
rect -4844 340718 -4608 340954
rect -5164 340398 -4928 340634
rect -4844 340398 -4608 340634
rect -5164 304718 -4928 304954
rect -4844 304718 -4608 304954
rect -5164 304398 -4928 304634
rect -4844 304398 -4608 304634
rect -5164 268718 -4928 268954
rect -4844 268718 -4608 268954
rect -5164 268398 -4928 268634
rect -4844 268398 -4608 268634
rect -5164 232718 -4928 232954
rect -4844 232718 -4608 232954
rect -5164 232398 -4928 232634
rect -4844 232398 -4608 232634
rect -5164 196718 -4928 196954
rect -4844 196718 -4608 196954
rect -5164 196398 -4928 196634
rect -4844 196398 -4608 196634
rect -5164 160718 -4928 160954
rect -4844 160718 -4608 160954
rect -5164 160398 -4928 160634
rect -4844 160398 -4608 160634
rect -5164 124718 -4928 124954
rect -4844 124718 -4608 124954
rect -5164 124398 -4928 124634
rect -4844 124398 -4608 124634
rect -5164 88718 -4928 88954
rect -4844 88718 -4608 88954
rect -5164 88398 -4928 88634
rect -4844 88398 -4608 88634
rect -5164 52718 -4928 52954
rect -4844 52718 -4608 52954
rect -5164 52398 -4928 52634
rect -4844 52398 -4608 52634
rect -5164 16718 -4928 16954
rect -4844 16718 -4608 16954
rect -5164 16398 -4928 16634
rect -4844 16398 -4608 16634
rect -4204 706832 -3968 707068
rect -3884 706832 -3648 707068
rect -4204 706512 -3968 706748
rect -3884 706512 -3648 706748
rect -4204 696218 -3968 696454
rect -3884 696218 -3648 696454
rect -4204 695898 -3968 696134
rect -3884 695898 -3648 696134
rect -4204 660218 -3968 660454
rect -3884 660218 -3648 660454
rect -4204 659898 -3968 660134
rect -3884 659898 -3648 660134
rect -4204 624218 -3968 624454
rect -3884 624218 -3648 624454
rect -4204 623898 -3968 624134
rect -3884 623898 -3648 624134
rect -4204 588218 -3968 588454
rect -3884 588218 -3648 588454
rect -4204 587898 -3968 588134
rect -3884 587898 -3648 588134
rect -4204 552218 -3968 552454
rect -3884 552218 -3648 552454
rect -4204 551898 -3968 552134
rect -3884 551898 -3648 552134
rect -4204 516218 -3968 516454
rect -3884 516218 -3648 516454
rect -4204 515898 -3968 516134
rect -3884 515898 -3648 516134
rect -4204 480218 -3968 480454
rect -3884 480218 -3648 480454
rect -4204 479898 -3968 480134
rect -3884 479898 -3648 480134
rect -4204 444218 -3968 444454
rect -3884 444218 -3648 444454
rect -4204 443898 -3968 444134
rect -3884 443898 -3648 444134
rect -4204 408218 -3968 408454
rect -3884 408218 -3648 408454
rect -4204 407898 -3968 408134
rect -3884 407898 -3648 408134
rect -4204 372218 -3968 372454
rect -3884 372218 -3648 372454
rect -4204 371898 -3968 372134
rect -3884 371898 -3648 372134
rect -4204 336218 -3968 336454
rect -3884 336218 -3648 336454
rect -4204 335898 -3968 336134
rect -3884 335898 -3648 336134
rect -4204 300218 -3968 300454
rect -3884 300218 -3648 300454
rect -4204 299898 -3968 300134
rect -3884 299898 -3648 300134
rect -4204 264218 -3968 264454
rect -3884 264218 -3648 264454
rect -4204 263898 -3968 264134
rect -3884 263898 -3648 264134
rect -4204 228218 -3968 228454
rect -3884 228218 -3648 228454
rect -4204 227898 -3968 228134
rect -3884 227898 -3648 228134
rect -4204 192218 -3968 192454
rect -3884 192218 -3648 192454
rect -4204 191898 -3968 192134
rect -3884 191898 -3648 192134
rect -4204 156218 -3968 156454
rect -3884 156218 -3648 156454
rect -4204 155898 -3968 156134
rect -3884 155898 -3648 156134
rect -4204 120218 -3968 120454
rect -3884 120218 -3648 120454
rect -4204 119898 -3968 120134
rect -3884 119898 -3648 120134
rect -4204 84218 -3968 84454
rect -3884 84218 -3648 84454
rect -4204 83898 -3968 84134
rect -3884 83898 -3648 84134
rect -4204 48218 -3968 48454
rect -3884 48218 -3648 48454
rect -4204 47898 -3968 48134
rect -3884 47898 -3648 48134
rect -4204 12218 -3968 12454
rect -3884 12218 -3648 12454
rect -4204 11898 -3968 12134
rect -3884 11898 -3648 12134
rect -3244 705872 -3008 706108
rect -2924 705872 -2688 706108
rect -3244 705552 -3008 705788
rect -2924 705552 -2688 705788
rect -3244 691718 -3008 691954
rect -2924 691718 -2688 691954
rect -3244 691398 -3008 691634
rect -2924 691398 -2688 691634
rect -3244 655718 -3008 655954
rect -2924 655718 -2688 655954
rect -3244 655398 -3008 655634
rect -2924 655398 -2688 655634
rect -3244 619718 -3008 619954
rect -2924 619718 -2688 619954
rect -3244 619398 -3008 619634
rect -2924 619398 -2688 619634
rect -3244 583718 -3008 583954
rect -2924 583718 -2688 583954
rect -3244 583398 -3008 583634
rect -2924 583398 -2688 583634
rect -3244 547718 -3008 547954
rect -2924 547718 -2688 547954
rect -3244 547398 -3008 547634
rect -2924 547398 -2688 547634
rect -3244 511718 -3008 511954
rect -2924 511718 -2688 511954
rect -3244 511398 -3008 511634
rect -2924 511398 -2688 511634
rect -3244 475718 -3008 475954
rect -2924 475718 -2688 475954
rect -3244 475398 -3008 475634
rect -2924 475398 -2688 475634
rect -3244 439718 -3008 439954
rect -2924 439718 -2688 439954
rect -3244 439398 -3008 439634
rect -2924 439398 -2688 439634
rect -3244 403718 -3008 403954
rect -2924 403718 -2688 403954
rect -3244 403398 -3008 403634
rect -2924 403398 -2688 403634
rect -3244 367718 -3008 367954
rect -2924 367718 -2688 367954
rect -3244 367398 -3008 367634
rect -2924 367398 -2688 367634
rect -3244 331718 -3008 331954
rect -2924 331718 -2688 331954
rect -3244 331398 -3008 331634
rect -2924 331398 -2688 331634
rect -3244 295718 -3008 295954
rect -2924 295718 -2688 295954
rect -3244 295398 -3008 295634
rect -2924 295398 -2688 295634
rect -3244 259718 -3008 259954
rect -2924 259718 -2688 259954
rect -3244 259398 -3008 259634
rect -2924 259398 -2688 259634
rect -3244 223718 -3008 223954
rect -2924 223718 -2688 223954
rect -3244 223398 -3008 223634
rect -2924 223398 -2688 223634
rect -3244 187718 -3008 187954
rect -2924 187718 -2688 187954
rect -3244 187398 -3008 187634
rect -2924 187398 -2688 187634
rect -3244 151718 -3008 151954
rect -2924 151718 -2688 151954
rect -3244 151398 -3008 151634
rect -2924 151398 -2688 151634
rect -3244 115718 -3008 115954
rect -2924 115718 -2688 115954
rect -3244 115398 -3008 115634
rect -2924 115398 -2688 115634
rect -3244 79718 -3008 79954
rect -2924 79718 -2688 79954
rect -3244 79398 -3008 79634
rect -2924 79398 -2688 79634
rect -3244 43718 -3008 43954
rect -2924 43718 -2688 43954
rect -3244 43398 -3008 43634
rect -2924 43398 -2688 43634
rect -3244 7718 -3008 7954
rect -2924 7718 -2688 7954
rect -3244 7398 -3008 7634
rect -2924 7398 -2688 7634
rect -2284 704912 -2048 705148
rect -1964 704912 -1728 705148
rect -2284 704592 -2048 704828
rect -1964 704592 -1728 704828
rect -2284 687218 -2048 687454
rect -1964 687218 -1728 687454
rect -2284 686898 -2048 687134
rect -1964 686898 -1728 687134
rect -2284 651218 -2048 651454
rect -1964 651218 -1728 651454
rect -2284 650898 -2048 651134
rect -1964 650898 -1728 651134
rect -2284 615218 -2048 615454
rect -1964 615218 -1728 615454
rect -2284 614898 -2048 615134
rect -1964 614898 -1728 615134
rect -2284 579218 -2048 579454
rect -1964 579218 -1728 579454
rect -2284 578898 -2048 579134
rect -1964 578898 -1728 579134
rect -2284 543218 -2048 543454
rect -1964 543218 -1728 543454
rect -2284 542898 -2048 543134
rect -1964 542898 -1728 543134
rect -2284 507218 -2048 507454
rect -1964 507218 -1728 507454
rect -2284 506898 -2048 507134
rect -1964 506898 -1728 507134
rect -2284 471218 -2048 471454
rect -1964 471218 -1728 471454
rect -2284 470898 -2048 471134
rect -1964 470898 -1728 471134
rect -2284 435218 -2048 435454
rect -1964 435218 -1728 435454
rect -2284 434898 -2048 435134
rect -1964 434898 -1728 435134
rect -2284 399218 -2048 399454
rect -1964 399218 -1728 399454
rect -2284 398898 -2048 399134
rect -1964 398898 -1728 399134
rect -2284 363218 -2048 363454
rect -1964 363218 -1728 363454
rect -2284 362898 -2048 363134
rect -1964 362898 -1728 363134
rect -2284 327218 -2048 327454
rect -1964 327218 -1728 327454
rect -2284 326898 -2048 327134
rect -1964 326898 -1728 327134
rect -2284 291218 -2048 291454
rect -1964 291218 -1728 291454
rect -2284 290898 -2048 291134
rect -1964 290898 -1728 291134
rect -2284 255218 -2048 255454
rect -1964 255218 -1728 255454
rect -2284 254898 -2048 255134
rect -1964 254898 -1728 255134
rect -2284 219218 -2048 219454
rect -1964 219218 -1728 219454
rect -2284 218898 -2048 219134
rect -1964 218898 -1728 219134
rect -2284 183218 -2048 183454
rect -1964 183218 -1728 183454
rect -2284 182898 -2048 183134
rect -1964 182898 -1728 183134
rect -2284 147218 -2048 147454
rect -1964 147218 -1728 147454
rect -2284 146898 -2048 147134
rect -1964 146898 -1728 147134
rect -2284 111218 -2048 111454
rect -1964 111218 -1728 111454
rect -2284 110898 -2048 111134
rect -1964 110898 -1728 111134
rect -2284 75218 -2048 75454
rect -1964 75218 -1728 75454
rect -2284 74898 -2048 75134
rect -1964 74898 -1728 75134
rect -2284 39218 -2048 39454
rect -1964 39218 -1728 39454
rect -2284 38898 -2048 39134
rect -1964 38898 -1728 39134
rect -2284 3218 -2048 3454
rect -1964 3218 -1728 3454
rect -2284 2898 -2048 3134
rect -1964 2898 -1728 3134
rect -2284 -892 -2048 -656
rect -1964 -892 -1728 -656
rect -2284 -1212 -2048 -976
rect -1964 -1212 -1728 -976
rect 1826 704912 2062 705148
rect 2146 704912 2382 705148
rect 1826 704592 2062 704828
rect 2146 704592 2382 704828
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -892 2062 -656
rect 2146 -892 2382 -656
rect 1826 -1212 2062 -976
rect 2146 -1212 2382 -976
rect -3244 -1852 -3008 -1616
rect -2924 -1852 -2688 -1616
rect -3244 -2172 -3008 -1936
rect -2924 -2172 -2688 -1936
rect -4204 -2812 -3968 -2576
rect -3884 -2812 -3648 -2576
rect -4204 -3132 -3968 -2896
rect -3884 -3132 -3648 -2896
rect -5164 -3772 -4928 -3536
rect -4844 -3772 -4608 -3536
rect -5164 -4092 -4928 -3856
rect -4844 -4092 -4608 -3856
rect -6124 -4732 -5888 -4496
rect -5804 -4732 -5568 -4496
rect -6124 -5052 -5888 -4816
rect -5804 -5052 -5568 -4816
rect -7084 -5692 -6848 -5456
rect -6764 -5692 -6528 -5456
rect -7084 -6012 -6848 -5776
rect -6764 -6012 -6528 -5776
rect -8044 -6652 -7808 -6416
rect -7724 -6652 -7488 -6416
rect -8044 -6972 -7808 -6736
rect -7724 -6972 -7488 -6736
rect -9004 -7612 -8768 -7376
rect -8684 -7612 -8448 -7376
rect -9004 -7932 -8768 -7696
rect -8684 -7932 -8448 -7696
rect 6326 705872 6562 706108
rect 6646 705872 6882 706108
rect 6326 705552 6562 705788
rect 6646 705552 6882 705788
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1852 6562 -1616
rect 6646 -1852 6882 -1616
rect 6326 -2172 6562 -1936
rect 6646 -2172 6882 -1936
rect 10826 706832 11062 707068
rect 11146 706832 11382 707068
rect 10826 706512 11062 706748
rect 11146 706512 11382 706748
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2812 11062 -2576
rect 11146 -2812 11382 -2576
rect 10826 -3132 11062 -2896
rect 11146 -3132 11382 -2896
rect 15326 707792 15562 708028
rect 15646 707792 15882 708028
rect 15326 707472 15562 707708
rect 15646 707472 15882 707708
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3772 15562 -3536
rect 15646 -3772 15882 -3536
rect 15326 -4092 15562 -3856
rect 15646 -4092 15882 -3856
rect 19826 708752 20062 708988
rect 20146 708752 20382 708988
rect 19826 708432 20062 708668
rect 20146 708432 20382 708668
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4732 20062 -4496
rect 20146 -4732 20382 -4496
rect 19826 -5052 20062 -4816
rect 20146 -5052 20382 -4816
rect 24326 709712 24562 709948
rect 24646 709712 24882 709948
rect 24326 709392 24562 709628
rect 24646 709392 24882 709628
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5692 24562 -5456
rect 24646 -5692 24882 -5456
rect 24326 -6012 24562 -5776
rect 24646 -6012 24882 -5776
rect 28826 710672 29062 710908
rect 29146 710672 29382 710908
rect 28826 710352 29062 710588
rect 29146 710352 29382 710588
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6652 29062 -6416
rect 29146 -6652 29382 -6416
rect 28826 -6972 29062 -6736
rect 29146 -6972 29382 -6736
rect 33326 711632 33562 711868
rect 33646 711632 33882 711868
rect 33326 711312 33562 711548
rect 33646 711312 33882 711548
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7612 33562 -7376
rect 33646 -7612 33882 -7376
rect 33326 -7932 33562 -7696
rect 33646 -7932 33882 -7696
rect 37826 704912 38062 705148
rect 38146 704912 38382 705148
rect 37826 704592 38062 704828
rect 38146 704592 38382 704828
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -892 38062 -656
rect 38146 -892 38382 -656
rect 37826 -1212 38062 -976
rect 38146 -1212 38382 -976
rect 42326 705872 42562 706108
rect 42646 705872 42882 706108
rect 42326 705552 42562 705788
rect 42646 705552 42882 705788
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1852 42562 -1616
rect 42646 -1852 42882 -1616
rect 42326 -2172 42562 -1936
rect 42646 -2172 42882 -1936
rect 46826 706832 47062 707068
rect 47146 706832 47382 707068
rect 46826 706512 47062 706748
rect 47146 706512 47382 706748
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2812 47062 -2576
rect 47146 -2812 47382 -2576
rect 46826 -3132 47062 -2896
rect 47146 -3132 47382 -2896
rect 51326 707792 51562 708028
rect 51646 707792 51882 708028
rect 51326 707472 51562 707708
rect 51646 707472 51882 707708
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3772 51562 -3536
rect 51646 -3772 51882 -3536
rect 51326 -4092 51562 -3856
rect 51646 -4092 51882 -3856
rect 55826 708752 56062 708988
rect 56146 708752 56382 708988
rect 55826 708432 56062 708668
rect 56146 708432 56382 708668
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4732 56062 -4496
rect 56146 -4732 56382 -4496
rect 55826 -5052 56062 -4816
rect 56146 -5052 56382 -4816
rect 60326 709712 60562 709948
rect 60646 709712 60882 709948
rect 60326 709392 60562 709628
rect 60646 709392 60882 709628
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5692 60562 -5456
rect 60646 -5692 60882 -5456
rect 60326 -6012 60562 -5776
rect 60646 -6012 60882 -5776
rect 64826 710672 65062 710908
rect 65146 710672 65382 710908
rect 64826 710352 65062 710588
rect 65146 710352 65382 710588
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6652 65062 -6416
rect 65146 -6652 65382 -6416
rect 64826 -6972 65062 -6736
rect 65146 -6972 65382 -6736
rect 69326 711632 69562 711868
rect 69646 711632 69882 711868
rect 69326 711312 69562 711548
rect 69646 711312 69882 711548
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7612 69562 -7376
rect 69646 -7612 69882 -7376
rect 69326 -7932 69562 -7696
rect 69646 -7932 69882 -7696
rect 73826 704912 74062 705148
rect 74146 704912 74382 705148
rect 73826 704592 74062 704828
rect 74146 704592 74382 704828
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -892 74062 -656
rect 74146 -892 74382 -656
rect 73826 -1212 74062 -976
rect 74146 -1212 74382 -976
rect 78326 705872 78562 706108
rect 78646 705872 78882 706108
rect 78326 705552 78562 705788
rect 78646 705552 78882 705788
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1852 78562 -1616
rect 78646 -1852 78882 -1616
rect 78326 -2172 78562 -1936
rect 78646 -2172 78882 -1936
rect 82826 706832 83062 707068
rect 83146 706832 83382 707068
rect 82826 706512 83062 706748
rect 83146 706512 83382 706748
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2812 83062 -2576
rect 83146 -2812 83382 -2576
rect 82826 -3132 83062 -2896
rect 83146 -3132 83382 -2896
rect 87326 707792 87562 708028
rect 87646 707792 87882 708028
rect 87326 707472 87562 707708
rect 87646 707472 87882 707708
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3772 87562 -3536
rect 87646 -3772 87882 -3536
rect 87326 -4092 87562 -3856
rect 87646 -4092 87882 -3856
rect 91826 708752 92062 708988
rect 92146 708752 92382 708988
rect 91826 708432 92062 708668
rect 92146 708432 92382 708668
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4732 92062 -4496
rect 92146 -4732 92382 -4496
rect 91826 -5052 92062 -4816
rect 92146 -5052 92382 -4816
rect 96326 709712 96562 709948
rect 96646 709712 96882 709948
rect 96326 709392 96562 709628
rect 96646 709392 96882 709628
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5692 96562 -5456
rect 96646 -5692 96882 -5456
rect 96326 -6012 96562 -5776
rect 96646 -6012 96882 -5776
rect 100826 710672 101062 710908
rect 101146 710672 101382 710908
rect 100826 710352 101062 710588
rect 101146 710352 101382 710588
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6652 101062 -6416
rect 101146 -6652 101382 -6416
rect 100826 -6972 101062 -6736
rect 101146 -6972 101382 -6736
rect 105326 711632 105562 711868
rect 105646 711632 105882 711868
rect 105326 711312 105562 711548
rect 105646 711312 105882 711548
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7612 105562 -7376
rect 105646 -7612 105882 -7376
rect 105326 -7932 105562 -7696
rect 105646 -7932 105882 -7696
rect 109826 704912 110062 705148
rect 110146 704912 110382 705148
rect 109826 704592 110062 704828
rect 110146 704592 110382 704828
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -892 110062 -656
rect 110146 -892 110382 -656
rect 109826 -1212 110062 -976
rect 110146 -1212 110382 -976
rect 114326 705872 114562 706108
rect 114646 705872 114882 706108
rect 114326 705552 114562 705788
rect 114646 705552 114882 705788
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1852 114562 -1616
rect 114646 -1852 114882 -1616
rect 114326 -2172 114562 -1936
rect 114646 -2172 114882 -1936
rect 118826 706832 119062 707068
rect 119146 706832 119382 707068
rect 118826 706512 119062 706748
rect 119146 706512 119382 706748
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2812 119062 -2576
rect 119146 -2812 119382 -2576
rect 118826 -3132 119062 -2896
rect 119146 -3132 119382 -2896
rect 123326 707792 123562 708028
rect 123646 707792 123882 708028
rect 123326 707472 123562 707708
rect 123646 707472 123882 707708
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3772 123562 -3536
rect 123646 -3772 123882 -3536
rect 123326 -4092 123562 -3856
rect 123646 -4092 123882 -3856
rect 127826 708752 128062 708988
rect 128146 708752 128382 708988
rect 127826 708432 128062 708668
rect 128146 708432 128382 708668
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4732 128062 -4496
rect 128146 -4732 128382 -4496
rect 127826 -5052 128062 -4816
rect 128146 -5052 128382 -4816
rect 132326 709712 132562 709948
rect 132646 709712 132882 709948
rect 132326 709392 132562 709628
rect 132646 709392 132882 709628
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5692 132562 -5456
rect 132646 -5692 132882 -5456
rect 132326 -6012 132562 -5776
rect 132646 -6012 132882 -5776
rect 136826 710672 137062 710908
rect 137146 710672 137382 710908
rect 136826 710352 137062 710588
rect 137146 710352 137382 710588
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6652 137062 -6416
rect 137146 -6652 137382 -6416
rect 136826 -6972 137062 -6736
rect 137146 -6972 137382 -6736
rect 141326 711632 141562 711868
rect 141646 711632 141882 711868
rect 141326 711312 141562 711548
rect 141646 711312 141882 711548
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7612 141562 -7376
rect 141646 -7612 141882 -7376
rect 141326 -7932 141562 -7696
rect 141646 -7932 141882 -7696
rect 145826 704912 146062 705148
rect 146146 704912 146382 705148
rect 145826 704592 146062 704828
rect 146146 704592 146382 704828
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -892 146062 -656
rect 146146 -892 146382 -656
rect 145826 -1212 146062 -976
rect 146146 -1212 146382 -976
rect 150326 705872 150562 706108
rect 150646 705872 150882 706108
rect 150326 705552 150562 705788
rect 150646 705552 150882 705788
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1852 150562 -1616
rect 150646 -1852 150882 -1616
rect 150326 -2172 150562 -1936
rect 150646 -2172 150882 -1936
rect 154826 706832 155062 707068
rect 155146 706832 155382 707068
rect 154826 706512 155062 706748
rect 155146 706512 155382 706748
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2812 155062 -2576
rect 155146 -2812 155382 -2576
rect 154826 -3132 155062 -2896
rect 155146 -3132 155382 -2896
rect 159326 707792 159562 708028
rect 159646 707792 159882 708028
rect 159326 707472 159562 707708
rect 159646 707472 159882 707708
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3772 159562 -3536
rect 159646 -3772 159882 -3536
rect 159326 -4092 159562 -3856
rect 159646 -4092 159882 -3856
rect 163826 708752 164062 708988
rect 164146 708752 164382 708988
rect 163826 708432 164062 708668
rect 164146 708432 164382 708668
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4732 164062 -4496
rect 164146 -4732 164382 -4496
rect 163826 -5052 164062 -4816
rect 164146 -5052 164382 -4816
rect 168326 709712 168562 709948
rect 168646 709712 168882 709948
rect 168326 709392 168562 709628
rect 168646 709392 168882 709628
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5692 168562 -5456
rect 168646 -5692 168882 -5456
rect 168326 -6012 168562 -5776
rect 168646 -6012 168882 -5776
rect 172826 710672 173062 710908
rect 173146 710672 173382 710908
rect 172826 710352 173062 710588
rect 173146 710352 173382 710588
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6652 173062 -6416
rect 173146 -6652 173382 -6416
rect 172826 -6972 173062 -6736
rect 173146 -6972 173382 -6736
rect 177326 711632 177562 711868
rect 177646 711632 177882 711868
rect 177326 711312 177562 711548
rect 177646 711312 177882 711548
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7612 177562 -7376
rect 177646 -7612 177882 -7376
rect 177326 -7932 177562 -7696
rect 177646 -7932 177882 -7696
rect 181826 704912 182062 705148
rect 182146 704912 182382 705148
rect 181826 704592 182062 704828
rect 182146 704592 182382 704828
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -892 182062 -656
rect 182146 -892 182382 -656
rect 181826 -1212 182062 -976
rect 182146 -1212 182382 -976
rect 186326 705872 186562 706108
rect 186646 705872 186882 706108
rect 186326 705552 186562 705788
rect 186646 705552 186882 705788
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1852 186562 -1616
rect 186646 -1852 186882 -1616
rect 186326 -2172 186562 -1936
rect 186646 -2172 186882 -1936
rect 190826 706832 191062 707068
rect 191146 706832 191382 707068
rect 190826 706512 191062 706748
rect 191146 706512 191382 706748
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2812 191062 -2576
rect 191146 -2812 191382 -2576
rect 190826 -3132 191062 -2896
rect 191146 -3132 191382 -2896
rect 195326 707792 195562 708028
rect 195646 707792 195882 708028
rect 195326 707472 195562 707708
rect 195646 707472 195882 707708
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3772 195562 -3536
rect 195646 -3772 195882 -3536
rect 195326 -4092 195562 -3856
rect 195646 -4092 195882 -3856
rect 199826 708752 200062 708988
rect 200146 708752 200382 708988
rect 199826 708432 200062 708668
rect 200146 708432 200382 708668
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4732 200062 -4496
rect 200146 -4732 200382 -4496
rect 199826 -5052 200062 -4816
rect 200146 -5052 200382 -4816
rect 204326 709712 204562 709948
rect 204646 709712 204882 709948
rect 204326 709392 204562 709628
rect 204646 709392 204882 709628
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5692 204562 -5456
rect 204646 -5692 204882 -5456
rect 204326 -6012 204562 -5776
rect 204646 -6012 204882 -5776
rect 208826 710672 209062 710908
rect 209146 710672 209382 710908
rect 208826 710352 209062 710588
rect 209146 710352 209382 710588
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6652 209062 -6416
rect 209146 -6652 209382 -6416
rect 208826 -6972 209062 -6736
rect 209146 -6972 209382 -6736
rect 213326 711632 213562 711868
rect 213646 711632 213882 711868
rect 213326 711312 213562 711548
rect 213646 711312 213882 711548
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7612 213562 -7376
rect 213646 -7612 213882 -7376
rect 213326 -7932 213562 -7696
rect 213646 -7932 213882 -7696
rect 217826 704912 218062 705148
rect 218146 704912 218382 705148
rect 217826 704592 218062 704828
rect 218146 704592 218382 704828
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -892 218062 -656
rect 218146 -892 218382 -656
rect 217826 -1212 218062 -976
rect 218146 -1212 218382 -976
rect 222326 705872 222562 706108
rect 222646 705872 222882 706108
rect 222326 705552 222562 705788
rect 222646 705552 222882 705788
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1852 222562 -1616
rect 222646 -1852 222882 -1616
rect 222326 -2172 222562 -1936
rect 222646 -2172 222882 -1936
rect 226826 706832 227062 707068
rect 227146 706832 227382 707068
rect 226826 706512 227062 706748
rect 227146 706512 227382 706748
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707792 231562 708028
rect 231646 707792 231882 708028
rect 231326 707472 231562 707708
rect 231646 707472 231882 707708
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708752 236062 708988
rect 236146 708752 236382 708988
rect 235826 708432 236062 708668
rect 236146 708432 236382 708668
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709712 240562 709948
rect 240646 709712 240882 709948
rect 240326 709392 240562 709628
rect 240646 709392 240882 709628
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710672 245062 710908
rect 245146 710672 245382 710908
rect 244826 710352 245062 710588
rect 245146 710352 245382 710588
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711632 249562 711868
rect 249646 711632 249882 711868
rect 249326 711312 249562 711548
rect 249646 711312 249882 711548
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 253826 704912 254062 705148
rect 254146 704912 254382 705148
rect 253826 704592 254062 704828
rect 254146 704592 254382 704828
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 258326 705872 258562 706108
rect 258646 705872 258882 706108
rect 258326 705552 258562 705788
rect 258646 705552 258882 705788
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 262826 706832 263062 707068
rect 263146 706832 263382 707068
rect 262826 706512 263062 706748
rect 263146 706512 263382 706748
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707792 267562 708028
rect 267646 707792 267882 708028
rect 267326 707472 267562 707708
rect 267646 707472 267882 707708
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708752 272062 708988
rect 272146 708752 272382 708988
rect 271826 708432 272062 708668
rect 272146 708432 272382 708668
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709712 276562 709948
rect 276646 709712 276882 709948
rect 276326 709392 276562 709628
rect 276646 709392 276882 709628
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710672 281062 710908
rect 281146 710672 281382 710908
rect 280826 710352 281062 710588
rect 281146 710352 281382 710588
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711632 285562 711868
rect 285646 711632 285882 711868
rect 285326 711312 285562 711548
rect 285646 711312 285882 711548
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 289826 704912 290062 705148
rect 290146 704912 290382 705148
rect 289826 704592 290062 704828
rect 290146 704592 290382 704828
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 294326 705872 294562 706108
rect 294646 705872 294882 706108
rect 294326 705552 294562 705788
rect 294646 705552 294882 705788
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 298826 706832 299062 707068
rect 299146 706832 299382 707068
rect 298826 706512 299062 706748
rect 299146 706512 299382 706748
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707792 303562 708028
rect 303646 707792 303882 708028
rect 303326 707472 303562 707708
rect 303646 707472 303882 707708
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708752 308062 708988
rect 308146 708752 308382 708988
rect 307826 708432 308062 708668
rect 308146 708432 308382 708668
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709712 312562 709948
rect 312646 709712 312882 709948
rect 312326 709392 312562 709628
rect 312646 709392 312882 709628
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710672 317062 710908
rect 317146 710672 317382 710908
rect 316826 710352 317062 710588
rect 317146 710352 317382 710588
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711632 321562 711868
rect 321646 711632 321882 711868
rect 321326 711312 321562 711548
rect 321646 711312 321882 711548
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 325826 704912 326062 705148
rect 326146 704912 326382 705148
rect 325826 704592 326062 704828
rect 326146 704592 326382 704828
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 330326 705872 330562 706108
rect 330646 705872 330882 706108
rect 330326 705552 330562 705788
rect 330646 705552 330882 705788
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 334826 706832 335062 707068
rect 335146 706832 335382 707068
rect 334826 706512 335062 706748
rect 335146 706512 335382 706748
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707792 339562 708028
rect 339646 707792 339882 708028
rect 339326 707472 339562 707708
rect 339646 707472 339882 707708
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708752 344062 708988
rect 344146 708752 344382 708988
rect 343826 708432 344062 708668
rect 344146 708432 344382 708668
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709712 348562 709948
rect 348646 709712 348882 709948
rect 348326 709392 348562 709628
rect 348646 709392 348882 709628
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710672 353062 710908
rect 353146 710672 353382 710908
rect 352826 710352 353062 710588
rect 353146 710352 353382 710588
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711632 357562 711868
rect 357646 711632 357882 711868
rect 357326 711312 357562 711548
rect 357646 711312 357882 711548
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 236250 255218 236486 255454
rect 236250 254898 236486 255134
rect 266970 255218 267206 255454
rect 266970 254898 267206 255134
rect 297690 255218 297926 255454
rect 297690 254898 297926 255134
rect 328410 255218 328646 255454
rect 328410 254898 328646 255134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 251610 223718 251846 223954
rect 251610 223398 251846 223634
rect 282330 223718 282566 223954
rect 282330 223398 282566 223634
rect 313050 223718 313286 223954
rect 313050 223398 313286 223634
rect 343770 223718 344006 223954
rect 343770 223398 344006 223634
rect 236250 219218 236486 219454
rect 236250 218898 236486 219134
rect 266970 219218 267206 219454
rect 266970 218898 267206 219134
rect 297690 219218 297926 219454
rect 297690 218898 297926 219134
rect 328410 219218 328646 219454
rect 328410 218898 328646 219134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 251610 187718 251846 187954
rect 251610 187398 251846 187634
rect 282330 187718 282566 187954
rect 282330 187398 282566 187634
rect 313050 187718 313286 187954
rect 313050 187398 313286 187634
rect 343770 187718 344006 187954
rect 343770 187398 344006 187634
rect 236250 183218 236486 183454
rect 236250 182898 236486 183134
rect 266970 183218 267206 183454
rect 266970 182898 267206 183134
rect 297690 183218 297926 183454
rect 297690 182898 297926 183134
rect 328410 183218 328646 183454
rect 328410 182898 328646 183134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 251610 151718 251846 151954
rect 251610 151398 251846 151634
rect 282330 151718 282566 151954
rect 282330 151398 282566 151634
rect 313050 151718 313286 151954
rect 313050 151398 313286 151634
rect 343770 151718 344006 151954
rect 343770 151398 344006 151634
rect 236250 147218 236486 147454
rect 236250 146898 236486 147134
rect 266970 147218 267206 147454
rect 266970 146898 267206 147134
rect 297690 147218 297926 147454
rect 297690 146898 297926 147134
rect 328410 147218 328646 147454
rect 328410 146898 328646 147134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 251610 115718 251846 115954
rect 251610 115398 251846 115634
rect 282330 115718 282566 115954
rect 282330 115398 282566 115634
rect 313050 115718 313286 115954
rect 313050 115398 313286 115634
rect 343770 115718 344006 115954
rect 343770 115398 344006 115634
rect 236250 111218 236486 111454
rect 236250 110898 236486 111134
rect 266970 111218 267206 111454
rect 266970 110898 267206 111134
rect 297690 111218 297926 111454
rect 297690 110898 297926 111134
rect 328410 111218 328646 111454
rect 328410 110898 328646 111134
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2812 227062 -2576
rect 227146 -2812 227382 -2576
rect 226826 -3132 227062 -2896
rect 227146 -3132 227382 -2896
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3772 231562 -3536
rect 231646 -3772 231882 -3536
rect 231326 -4092 231562 -3856
rect 231646 -4092 231882 -3856
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4732 236062 -4496
rect 236146 -4732 236382 -4496
rect 235826 -5052 236062 -4816
rect 236146 -5052 236382 -4816
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5692 240562 -5456
rect 240646 -5692 240882 -5456
rect 240326 -6012 240562 -5776
rect 240646 -6012 240882 -5776
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6652 245062 -6416
rect 245146 -6652 245382 -6416
rect 244826 -6972 245062 -6736
rect 245146 -6972 245382 -6736
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7612 249562 -7376
rect 249646 -7612 249882 -7376
rect 249326 -7932 249562 -7696
rect 249646 -7932 249882 -7696
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -892 254062 -656
rect 254146 -892 254382 -656
rect 253826 -1212 254062 -976
rect 254146 -1212 254382 -976
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1852 258562 -1616
rect 258646 -1852 258882 -1616
rect 258326 -2172 258562 -1936
rect 258646 -2172 258882 -1936
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2812 263062 -2576
rect 263146 -2812 263382 -2576
rect 262826 -3132 263062 -2896
rect 263146 -3132 263382 -2896
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3772 267562 -3536
rect 267646 -3772 267882 -3536
rect 267326 -4092 267562 -3856
rect 267646 -4092 267882 -3856
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4732 272062 -4496
rect 272146 -4732 272382 -4496
rect 271826 -5052 272062 -4816
rect 272146 -5052 272382 -4816
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5692 276562 -5456
rect 276646 -5692 276882 -5456
rect 276326 -6012 276562 -5776
rect 276646 -6012 276882 -5776
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6652 281062 -6416
rect 281146 -6652 281382 -6416
rect 280826 -6972 281062 -6736
rect 281146 -6972 281382 -6736
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7612 285562 -7376
rect 285646 -7612 285882 -7376
rect 285326 -7932 285562 -7696
rect 285646 -7932 285882 -7696
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -892 290062 -656
rect 290146 -892 290382 -656
rect 289826 -1212 290062 -976
rect 290146 -1212 290382 -976
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1852 294562 -1616
rect 294646 -1852 294882 -1616
rect 294326 -2172 294562 -1936
rect 294646 -2172 294882 -1936
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2812 299062 -2576
rect 299146 -2812 299382 -2576
rect 298826 -3132 299062 -2896
rect 299146 -3132 299382 -2896
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3772 303562 -3536
rect 303646 -3772 303882 -3536
rect 303326 -4092 303562 -3856
rect 303646 -4092 303882 -3856
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4732 308062 -4496
rect 308146 -4732 308382 -4496
rect 307826 -5052 308062 -4816
rect 308146 -5052 308382 -4816
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5692 312562 -5456
rect 312646 -5692 312882 -5456
rect 312326 -6012 312562 -5776
rect 312646 -6012 312882 -5776
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6652 317062 -6416
rect 317146 -6652 317382 -6416
rect 316826 -6972 317062 -6736
rect 317146 -6972 317382 -6736
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7612 321562 -7376
rect 321646 -7612 321882 -7376
rect 321326 -7932 321562 -7696
rect 321646 -7932 321882 -7696
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -892 326062 -656
rect 326146 -892 326382 -656
rect 325826 -1212 326062 -976
rect 326146 -1212 326382 -976
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1852 330562 -1616
rect 330646 -1852 330882 -1616
rect 330326 -2172 330562 -1936
rect 330646 -2172 330882 -1936
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2812 335062 -2576
rect 335146 -2812 335382 -2576
rect 334826 -3132 335062 -2896
rect 335146 -3132 335382 -2896
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3772 339562 -3536
rect 339646 -3772 339882 -3536
rect 339326 -4092 339562 -3856
rect 339646 -4092 339882 -3856
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4732 344062 -4496
rect 344146 -4732 344382 -4496
rect 343826 -5052 344062 -4816
rect 344146 -5052 344382 -4816
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5692 348562 -5456
rect 348646 -5692 348882 -5456
rect 348326 -6012 348562 -5776
rect 348646 -6012 348882 -5776
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6652 353062 -6416
rect 353146 -6652 353382 -6416
rect 352826 -6972 353062 -6736
rect 353146 -6972 353382 -6736
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7612 357562 -7376
rect 357646 -7612 357882 -7376
rect 357326 -7932 357562 -7696
rect 357646 -7932 357882 -7696
rect 361826 704912 362062 705148
rect 362146 704912 362382 705148
rect 361826 704592 362062 704828
rect 362146 704592 362382 704828
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -892 362062 -656
rect 362146 -892 362382 -656
rect 361826 -1212 362062 -976
rect 362146 -1212 362382 -976
rect 366326 705872 366562 706108
rect 366646 705872 366882 706108
rect 366326 705552 366562 705788
rect 366646 705552 366882 705788
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1852 366562 -1616
rect 366646 -1852 366882 -1616
rect 366326 -2172 366562 -1936
rect 366646 -2172 366882 -1936
rect 370826 706832 371062 707068
rect 371146 706832 371382 707068
rect 370826 706512 371062 706748
rect 371146 706512 371382 706748
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2812 371062 -2576
rect 371146 -2812 371382 -2576
rect 370826 -3132 371062 -2896
rect 371146 -3132 371382 -2896
rect 375326 707792 375562 708028
rect 375646 707792 375882 708028
rect 375326 707472 375562 707708
rect 375646 707472 375882 707708
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3772 375562 -3536
rect 375646 -3772 375882 -3536
rect 375326 -4092 375562 -3856
rect 375646 -4092 375882 -3856
rect 379826 708752 380062 708988
rect 380146 708752 380382 708988
rect 379826 708432 380062 708668
rect 380146 708432 380382 708668
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4732 380062 -4496
rect 380146 -4732 380382 -4496
rect 379826 -5052 380062 -4816
rect 380146 -5052 380382 -4816
rect 384326 709712 384562 709948
rect 384646 709712 384882 709948
rect 384326 709392 384562 709628
rect 384646 709392 384882 709628
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5692 384562 -5456
rect 384646 -5692 384882 -5456
rect 384326 -6012 384562 -5776
rect 384646 -6012 384882 -5776
rect 388826 710672 389062 710908
rect 389146 710672 389382 710908
rect 388826 710352 389062 710588
rect 389146 710352 389382 710588
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6652 389062 -6416
rect 389146 -6652 389382 -6416
rect 388826 -6972 389062 -6736
rect 389146 -6972 389382 -6736
rect 393326 711632 393562 711868
rect 393646 711632 393882 711868
rect 393326 711312 393562 711548
rect 393646 711312 393882 711548
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7612 393562 -7376
rect 393646 -7612 393882 -7376
rect 393326 -7932 393562 -7696
rect 393646 -7932 393882 -7696
rect 397826 704912 398062 705148
rect 398146 704912 398382 705148
rect 397826 704592 398062 704828
rect 398146 704592 398382 704828
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -892 398062 -656
rect 398146 -892 398382 -656
rect 397826 -1212 398062 -976
rect 398146 -1212 398382 -976
rect 402326 705872 402562 706108
rect 402646 705872 402882 706108
rect 402326 705552 402562 705788
rect 402646 705552 402882 705788
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1852 402562 -1616
rect 402646 -1852 402882 -1616
rect 402326 -2172 402562 -1936
rect 402646 -2172 402882 -1936
rect 406826 706832 407062 707068
rect 407146 706832 407382 707068
rect 406826 706512 407062 706748
rect 407146 706512 407382 706748
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2812 407062 -2576
rect 407146 -2812 407382 -2576
rect 406826 -3132 407062 -2896
rect 407146 -3132 407382 -2896
rect 411326 707792 411562 708028
rect 411646 707792 411882 708028
rect 411326 707472 411562 707708
rect 411646 707472 411882 707708
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3772 411562 -3536
rect 411646 -3772 411882 -3536
rect 411326 -4092 411562 -3856
rect 411646 -4092 411882 -3856
rect 415826 708752 416062 708988
rect 416146 708752 416382 708988
rect 415826 708432 416062 708668
rect 416146 708432 416382 708668
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4732 416062 -4496
rect 416146 -4732 416382 -4496
rect 415826 -5052 416062 -4816
rect 416146 -5052 416382 -4816
rect 420326 709712 420562 709948
rect 420646 709712 420882 709948
rect 420326 709392 420562 709628
rect 420646 709392 420882 709628
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5692 420562 -5456
rect 420646 -5692 420882 -5456
rect 420326 -6012 420562 -5776
rect 420646 -6012 420882 -5776
rect 424826 710672 425062 710908
rect 425146 710672 425382 710908
rect 424826 710352 425062 710588
rect 425146 710352 425382 710588
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6652 425062 -6416
rect 425146 -6652 425382 -6416
rect 424826 -6972 425062 -6736
rect 425146 -6972 425382 -6736
rect 429326 711632 429562 711868
rect 429646 711632 429882 711868
rect 429326 711312 429562 711548
rect 429646 711312 429882 711548
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7612 429562 -7376
rect 429646 -7612 429882 -7376
rect 429326 -7932 429562 -7696
rect 429646 -7932 429882 -7696
rect 433826 704912 434062 705148
rect 434146 704912 434382 705148
rect 433826 704592 434062 704828
rect 434146 704592 434382 704828
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -892 434062 -656
rect 434146 -892 434382 -656
rect 433826 -1212 434062 -976
rect 434146 -1212 434382 -976
rect 438326 705872 438562 706108
rect 438646 705872 438882 706108
rect 438326 705552 438562 705788
rect 438646 705552 438882 705788
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1852 438562 -1616
rect 438646 -1852 438882 -1616
rect 438326 -2172 438562 -1936
rect 438646 -2172 438882 -1936
rect 442826 706832 443062 707068
rect 443146 706832 443382 707068
rect 442826 706512 443062 706748
rect 443146 706512 443382 706748
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2812 443062 -2576
rect 443146 -2812 443382 -2576
rect 442826 -3132 443062 -2896
rect 443146 -3132 443382 -2896
rect 447326 707792 447562 708028
rect 447646 707792 447882 708028
rect 447326 707472 447562 707708
rect 447646 707472 447882 707708
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3772 447562 -3536
rect 447646 -3772 447882 -3536
rect 447326 -4092 447562 -3856
rect 447646 -4092 447882 -3856
rect 451826 708752 452062 708988
rect 452146 708752 452382 708988
rect 451826 708432 452062 708668
rect 452146 708432 452382 708668
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4732 452062 -4496
rect 452146 -4732 452382 -4496
rect 451826 -5052 452062 -4816
rect 452146 -5052 452382 -4816
rect 456326 709712 456562 709948
rect 456646 709712 456882 709948
rect 456326 709392 456562 709628
rect 456646 709392 456882 709628
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5692 456562 -5456
rect 456646 -5692 456882 -5456
rect 456326 -6012 456562 -5776
rect 456646 -6012 456882 -5776
rect 460826 710672 461062 710908
rect 461146 710672 461382 710908
rect 460826 710352 461062 710588
rect 461146 710352 461382 710588
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6652 461062 -6416
rect 461146 -6652 461382 -6416
rect 460826 -6972 461062 -6736
rect 461146 -6972 461382 -6736
rect 465326 711632 465562 711868
rect 465646 711632 465882 711868
rect 465326 711312 465562 711548
rect 465646 711312 465882 711548
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7612 465562 -7376
rect 465646 -7612 465882 -7376
rect 465326 -7932 465562 -7696
rect 465646 -7932 465882 -7696
rect 469826 704912 470062 705148
rect 470146 704912 470382 705148
rect 469826 704592 470062 704828
rect 470146 704592 470382 704828
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -892 470062 -656
rect 470146 -892 470382 -656
rect 469826 -1212 470062 -976
rect 470146 -1212 470382 -976
rect 474326 705872 474562 706108
rect 474646 705872 474882 706108
rect 474326 705552 474562 705788
rect 474646 705552 474882 705788
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1852 474562 -1616
rect 474646 -1852 474882 -1616
rect 474326 -2172 474562 -1936
rect 474646 -2172 474882 -1936
rect 478826 706832 479062 707068
rect 479146 706832 479382 707068
rect 478826 706512 479062 706748
rect 479146 706512 479382 706748
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2812 479062 -2576
rect 479146 -2812 479382 -2576
rect 478826 -3132 479062 -2896
rect 479146 -3132 479382 -2896
rect 483326 707792 483562 708028
rect 483646 707792 483882 708028
rect 483326 707472 483562 707708
rect 483646 707472 483882 707708
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3772 483562 -3536
rect 483646 -3772 483882 -3536
rect 483326 -4092 483562 -3856
rect 483646 -4092 483882 -3856
rect 487826 708752 488062 708988
rect 488146 708752 488382 708988
rect 487826 708432 488062 708668
rect 488146 708432 488382 708668
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4732 488062 -4496
rect 488146 -4732 488382 -4496
rect 487826 -5052 488062 -4816
rect 488146 -5052 488382 -4816
rect 492326 709712 492562 709948
rect 492646 709712 492882 709948
rect 492326 709392 492562 709628
rect 492646 709392 492882 709628
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5692 492562 -5456
rect 492646 -5692 492882 -5456
rect 492326 -6012 492562 -5776
rect 492646 -6012 492882 -5776
rect 496826 710672 497062 710908
rect 497146 710672 497382 710908
rect 496826 710352 497062 710588
rect 497146 710352 497382 710588
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6652 497062 -6416
rect 497146 -6652 497382 -6416
rect 496826 -6972 497062 -6736
rect 497146 -6972 497382 -6736
rect 501326 711632 501562 711868
rect 501646 711632 501882 711868
rect 501326 711312 501562 711548
rect 501646 711312 501882 711548
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7612 501562 -7376
rect 501646 -7612 501882 -7376
rect 501326 -7932 501562 -7696
rect 501646 -7932 501882 -7696
rect 505826 704912 506062 705148
rect 506146 704912 506382 705148
rect 505826 704592 506062 704828
rect 506146 704592 506382 704828
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -892 506062 -656
rect 506146 -892 506382 -656
rect 505826 -1212 506062 -976
rect 506146 -1212 506382 -976
rect 510326 705872 510562 706108
rect 510646 705872 510882 706108
rect 510326 705552 510562 705788
rect 510646 705552 510882 705788
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1852 510562 -1616
rect 510646 -1852 510882 -1616
rect 510326 -2172 510562 -1936
rect 510646 -2172 510882 -1936
rect 514826 706832 515062 707068
rect 515146 706832 515382 707068
rect 514826 706512 515062 706748
rect 515146 706512 515382 706748
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2812 515062 -2576
rect 515146 -2812 515382 -2576
rect 514826 -3132 515062 -2896
rect 515146 -3132 515382 -2896
rect 519326 707792 519562 708028
rect 519646 707792 519882 708028
rect 519326 707472 519562 707708
rect 519646 707472 519882 707708
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3772 519562 -3536
rect 519646 -3772 519882 -3536
rect 519326 -4092 519562 -3856
rect 519646 -4092 519882 -3856
rect 523826 708752 524062 708988
rect 524146 708752 524382 708988
rect 523826 708432 524062 708668
rect 524146 708432 524382 708668
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4732 524062 -4496
rect 524146 -4732 524382 -4496
rect 523826 -5052 524062 -4816
rect 524146 -5052 524382 -4816
rect 528326 709712 528562 709948
rect 528646 709712 528882 709948
rect 528326 709392 528562 709628
rect 528646 709392 528882 709628
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5692 528562 -5456
rect 528646 -5692 528882 -5456
rect 528326 -6012 528562 -5776
rect 528646 -6012 528882 -5776
rect 532826 710672 533062 710908
rect 533146 710672 533382 710908
rect 532826 710352 533062 710588
rect 533146 710352 533382 710588
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6652 533062 -6416
rect 533146 -6652 533382 -6416
rect 532826 -6972 533062 -6736
rect 533146 -6972 533382 -6736
rect 537326 711632 537562 711868
rect 537646 711632 537882 711868
rect 537326 711312 537562 711548
rect 537646 711312 537882 711548
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7612 537562 -7376
rect 537646 -7612 537882 -7376
rect 537326 -7932 537562 -7696
rect 537646 -7932 537882 -7696
rect 541826 704912 542062 705148
rect 542146 704912 542382 705148
rect 541826 704592 542062 704828
rect 542146 704592 542382 704828
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -892 542062 -656
rect 542146 -892 542382 -656
rect 541826 -1212 542062 -976
rect 542146 -1212 542382 -976
rect 546326 705872 546562 706108
rect 546646 705872 546882 706108
rect 546326 705552 546562 705788
rect 546646 705552 546882 705788
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1852 546562 -1616
rect 546646 -1852 546882 -1616
rect 546326 -2172 546562 -1936
rect 546646 -2172 546882 -1936
rect 550826 706832 551062 707068
rect 551146 706832 551382 707068
rect 550826 706512 551062 706748
rect 551146 706512 551382 706748
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2812 551062 -2576
rect 551146 -2812 551382 -2576
rect 550826 -3132 551062 -2896
rect 551146 -3132 551382 -2896
rect 555326 707792 555562 708028
rect 555646 707792 555882 708028
rect 555326 707472 555562 707708
rect 555646 707472 555882 707708
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3772 555562 -3536
rect 555646 -3772 555882 -3536
rect 555326 -4092 555562 -3856
rect 555646 -4092 555882 -3856
rect 559826 708752 560062 708988
rect 560146 708752 560382 708988
rect 559826 708432 560062 708668
rect 560146 708432 560382 708668
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4732 560062 -4496
rect 560146 -4732 560382 -4496
rect 559826 -5052 560062 -4816
rect 560146 -5052 560382 -4816
rect 564326 709712 564562 709948
rect 564646 709712 564882 709948
rect 564326 709392 564562 709628
rect 564646 709392 564882 709628
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5692 564562 -5456
rect 564646 -5692 564882 -5456
rect 564326 -6012 564562 -5776
rect 564646 -6012 564882 -5776
rect 568826 710672 569062 710908
rect 569146 710672 569382 710908
rect 568826 710352 569062 710588
rect 569146 710352 569382 710588
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6652 569062 -6416
rect 569146 -6652 569382 -6416
rect 568826 -6972 569062 -6736
rect 569146 -6972 569382 -6736
rect 573326 711632 573562 711868
rect 573646 711632 573882 711868
rect 573326 711312 573562 711548
rect 573646 711312 573882 711548
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7612 573562 -7376
rect 573646 -7612 573882 -7376
rect 573326 -7932 573562 -7696
rect 573646 -7932 573882 -7696
rect 577826 704912 578062 705148
rect 578146 704912 578382 705148
rect 577826 704592 578062 704828
rect 578146 704592 578382 704828
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -892 578062 -656
rect 578146 -892 578382 -656
rect 577826 -1212 578062 -976
rect 578146 -1212 578382 -976
rect 592372 711632 592608 711868
rect 592692 711632 592928 711868
rect 592372 711312 592608 711548
rect 592692 711312 592928 711548
rect 591412 710672 591648 710908
rect 591732 710672 591968 710908
rect 591412 710352 591648 710588
rect 591732 710352 591968 710588
rect 590452 709712 590688 709948
rect 590772 709712 591008 709948
rect 590452 709392 590688 709628
rect 590772 709392 591008 709628
rect 589492 708752 589728 708988
rect 589812 708752 590048 708988
rect 589492 708432 589728 708668
rect 589812 708432 590048 708668
rect 588532 707792 588768 708028
rect 588852 707792 589088 708028
rect 588532 707472 588768 707708
rect 588852 707472 589088 707708
rect 587572 706832 587808 707068
rect 587892 706832 588128 707068
rect 587572 706512 587808 706748
rect 587892 706512 588128 706748
rect 582326 705872 582562 706108
rect 582646 705872 582882 706108
rect 582326 705552 582562 705788
rect 582646 705552 582882 705788
rect 586612 705872 586848 706108
rect 586932 705872 587168 706108
rect 586612 705552 586848 705788
rect 586932 705552 587168 705788
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585652 704912 585888 705148
rect 585972 704912 586208 705148
rect 585652 704592 585888 704828
rect 585972 704592 586208 704828
rect 585652 687218 585888 687454
rect 585972 687218 586208 687454
rect 585652 686898 585888 687134
rect 585972 686898 586208 687134
rect 585652 651218 585888 651454
rect 585972 651218 586208 651454
rect 585652 650898 585888 651134
rect 585972 650898 586208 651134
rect 585652 615218 585888 615454
rect 585972 615218 586208 615454
rect 585652 614898 585888 615134
rect 585972 614898 586208 615134
rect 585652 579218 585888 579454
rect 585972 579218 586208 579454
rect 585652 578898 585888 579134
rect 585972 578898 586208 579134
rect 585652 543218 585888 543454
rect 585972 543218 586208 543454
rect 585652 542898 585888 543134
rect 585972 542898 586208 543134
rect 585652 507218 585888 507454
rect 585972 507218 586208 507454
rect 585652 506898 585888 507134
rect 585972 506898 586208 507134
rect 585652 471218 585888 471454
rect 585972 471218 586208 471454
rect 585652 470898 585888 471134
rect 585972 470898 586208 471134
rect 585652 435218 585888 435454
rect 585972 435218 586208 435454
rect 585652 434898 585888 435134
rect 585972 434898 586208 435134
rect 585652 399218 585888 399454
rect 585972 399218 586208 399454
rect 585652 398898 585888 399134
rect 585972 398898 586208 399134
rect 585652 363218 585888 363454
rect 585972 363218 586208 363454
rect 585652 362898 585888 363134
rect 585972 362898 586208 363134
rect 585652 327218 585888 327454
rect 585972 327218 586208 327454
rect 585652 326898 585888 327134
rect 585972 326898 586208 327134
rect 585652 291218 585888 291454
rect 585972 291218 586208 291454
rect 585652 290898 585888 291134
rect 585972 290898 586208 291134
rect 585652 255218 585888 255454
rect 585972 255218 586208 255454
rect 585652 254898 585888 255134
rect 585972 254898 586208 255134
rect 585652 219218 585888 219454
rect 585972 219218 586208 219454
rect 585652 218898 585888 219134
rect 585972 218898 586208 219134
rect 585652 183218 585888 183454
rect 585972 183218 586208 183454
rect 585652 182898 585888 183134
rect 585972 182898 586208 183134
rect 585652 147218 585888 147454
rect 585972 147218 586208 147454
rect 585652 146898 585888 147134
rect 585972 146898 586208 147134
rect 585652 111218 585888 111454
rect 585972 111218 586208 111454
rect 585652 110898 585888 111134
rect 585972 110898 586208 111134
rect 585652 75218 585888 75454
rect 585972 75218 586208 75454
rect 585652 74898 585888 75134
rect 585972 74898 586208 75134
rect 585652 39218 585888 39454
rect 585972 39218 586208 39454
rect 585652 38898 585888 39134
rect 585972 38898 586208 39134
rect 585652 3218 585888 3454
rect 585972 3218 586208 3454
rect 585652 2898 585888 3134
rect 585972 2898 586208 3134
rect 585652 -892 585888 -656
rect 585972 -892 586208 -656
rect 585652 -1212 585888 -976
rect 585972 -1212 586208 -976
rect 586612 691718 586848 691954
rect 586932 691718 587168 691954
rect 586612 691398 586848 691634
rect 586932 691398 587168 691634
rect 586612 655718 586848 655954
rect 586932 655718 587168 655954
rect 586612 655398 586848 655634
rect 586932 655398 587168 655634
rect 586612 619718 586848 619954
rect 586932 619718 587168 619954
rect 586612 619398 586848 619634
rect 586932 619398 587168 619634
rect 586612 583718 586848 583954
rect 586932 583718 587168 583954
rect 586612 583398 586848 583634
rect 586932 583398 587168 583634
rect 586612 547718 586848 547954
rect 586932 547718 587168 547954
rect 586612 547398 586848 547634
rect 586932 547398 587168 547634
rect 586612 511718 586848 511954
rect 586932 511718 587168 511954
rect 586612 511398 586848 511634
rect 586932 511398 587168 511634
rect 586612 475718 586848 475954
rect 586932 475718 587168 475954
rect 586612 475398 586848 475634
rect 586932 475398 587168 475634
rect 586612 439718 586848 439954
rect 586932 439718 587168 439954
rect 586612 439398 586848 439634
rect 586932 439398 587168 439634
rect 586612 403718 586848 403954
rect 586932 403718 587168 403954
rect 586612 403398 586848 403634
rect 586932 403398 587168 403634
rect 586612 367718 586848 367954
rect 586932 367718 587168 367954
rect 586612 367398 586848 367634
rect 586932 367398 587168 367634
rect 586612 331718 586848 331954
rect 586932 331718 587168 331954
rect 586612 331398 586848 331634
rect 586932 331398 587168 331634
rect 586612 295718 586848 295954
rect 586932 295718 587168 295954
rect 586612 295398 586848 295634
rect 586932 295398 587168 295634
rect 586612 259718 586848 259954
rect 586932 259718 587168 259954
rect 586612 259398 586848 259634
rect 586932 259398 587168 259634
rect 586612 223718 586848 223954
rect 586932 223718 587168 223954
rect 586612 223398 586848 223634
rect 586932 223398 587168 223634
rect 586612 187718 586848 187954
rect 586932 187718 587168 187954
rect 586612 187398 586848 187634
rect 586932 187398 587168 187634
rect 586612 151718 586848 151954
rect 586932 151718 587168 151954
rect 586612 151398 586848 151634
rect 586932 151398 587168 151634
rect 586612 115718 586848 115954
rect 586932 115718 587168 115954
rect 586612 115398 586848 115634
rect 586932 115398 587168 115634
rect 586612 79718 586848 79954
rect 586932 79718 587168 79954
rect 586612 79398 586848 79634
rect 586932 79398 587168 79634
rect 586612 43718 586848 43954
rect 586932 43718 587168 43954
rect 586612 43398 586848 43634
rect 586932 43398 587168 43634
rect 586612 7718 586848 7954
rect 586932 7718 587168 7954
rect 586612 7398 586848 7634
rect 586932 7398 587168 7634
rect 582326 -1852 582562 -1616
rect 582646 -1852 582882 -1616
rect 582326 -2172 582562 -1936
rect 582646 -2172 582882 -1936
rect 586612 -1852 586848 -1616
rect 586932 -1852 587168 -1616
rect 586612 -2172 586848 -1936
rect 586932 -2172 587168 -1936
rect 587572 696218 587808 696454
rect 587892 696218 588128 696454
rect 587572 695898 587808 696134
rect 587892 695898 588128 696134
rect 587572 660218 587808 660454
rect 587892 660218 588128 660454
rect 587572 659898 587808 660134
rect 587892 659898 588128 660134
rect 587572 624218 587808 624454
rect 587892 624218 588128 624454
rect 587572 623898 587808 624134
rect 587892 623898 588128 624134
rect 587572 588218 587808 588454
rect 587892 588218 588128 588454
rect 587572 587898 587808 588134
rect 587892 587898 588128 588134
rect 587572 552218 587808 552454
rect 587892 552218 588128 552454
rect 587572 551898 587808 552134
rect 587892 551898 588128 552134
rect 587572 516218 587808 516454
rect 587892 516218 588128 516454
rect 587572 515898 587808 516134
rect 587892 515898 588128 516134
rect 587572 480218 587808 480454
rect 587892 480218 588128 480454
rect 587572 479898 587808 480134
rect 587892 479898 588128 480134
rect 587572 444218 587808 444454
rect 587892 444218 588128 444454
rect 587572 443898 587808 444134
rect 587892 443898 588128 444134
rect 587572 408218 587808 408454
rect 587892 408218 588128 408454
rect 587572 407898 587808 408134
rect 587892 407898 588128 408134
rect 587572 372218 587808 372454
rect 587892 372218 588128 372454
rect 587572 371898 587808 372134
rect 587892 371898 588128 372134
rect 587572 336218 587808 336454
rect 587892 336218 588128 336454
rect 587572 335898 587808 336134
rect 587892 335898 588128 336134
rect 587572 300218 587808 300454
rect 587892 300218 588128 300454
rect 587572 299898 587808 300134
rect 587892 299898 588128 300134
rect 587572 264218 587808 264454
rect 587892 264218 588128 264454
rect 587572 263898 587808 264134
rect 587892 263898 588128 264134
rect 587572 228218 587808 228454
rect 587892 228218 588128 228454
rect 587572 227898 587808 228134
rect 587892 227898 588128 228134
rect 587572 192218 587808 192454
rect 587892 192218 588128 192454
rect 587572 191898 587808 192134
rect 587892 191898 588128 192134
rect 587572 156218 587808 156454
rect 587892 156218 588128 156454
rect 587572 155898 587808 156134
rect 587892 155898 588128 156134
rect 587572 120218 587808 120454
rect 587892 120218 588128 120454
rect 587572 119898 587808 120134
rect 587892 119898 588128 120134
rect 587572 84218 587808 84454
rect 587892 84218 588128 84454
rect 587572 83898 587808 84134
rect 587892 83898 588128 84134
rect 587572 48218 587808 48454
rect 587892 48218 588128 48454
rect 587572 47898 587808 48134
rect 587892 47898 588128 48134
rect 587572 12218 587808 12454
rect 587892 12218 588128 12454
rect 587572 11898 587808 12134
rect 587892 11898 588128 12134
rect 587572 -2812 587808 -2576
rect 587892 -2812 588128 -2576
rect 587572 -3132 587808 -2896
rect 587892 -3132 588128 -2896
rect 588532 700718 588768 700954
rect 588852 700718 589088 700954
rect 588532 700398 588768 700634
rect 588852 700398 589088 700634
rect 588532 664718 588768 664954
rect 588852 664718 589088 664954
rect 588532 664398 588768 664634
rect 588852 664398 589088 664634
rect 588532 628718 588768 628954
rect 588852 628718 589088 628954
rect 588532 628398 588768 628634
rect 588852 628398 589088 628634
rect 588532 592718 588768 592954
rect 588852 592718 589088 592954
rect 588532 592398 588768 592634
rect 588852 592398 589088 592634
rect 588532 556718 588768 556954
rect 588852 556718 589088 556954
rect 588532 556398 588768 556634
rect 588852 556398 589088 556634
rect 588532 520718 588768 520954
rect 588852 520718 589088 520954
rect 588532 520398 588768 520634
rect 588852 520398 589088 520634
rect 588532 484718 588768 484954
rect 588852 484718 589088 484954
rect 588532 484398 588768 484634
rect 588852 484398 589088 484634
rect 588532 448718 588768 448954
rect 588852 448718 589088 448954
rect 588532 448398 588768 448634
rect 588852 448398 589088 448634
rect 588532 412718 588768 412954
rect 588852 412718 589088 412954
rect 588532 412398 588768 412634
rect 588852 412398 589088 412634
rect 588532 376718 588768 376954
rect 588852 376718 589088 376954
rect 588532 376398 588768 376634
rect 588852 376398 589088 376634
rect 588532 340718 588768 340954
rect 588852 340718 589088 340954
rect 588532 340398 588768 340634
rect 588852 340398 589088 340634
rect 588532 304718 588768 304954
rect 588852 304718 589088 304954
rect 588532 304398 588768 304634
rect 588852 304398 589088 304634
rect 588532 268718 588768 268954
rect 588852 268718 589088 268954
rect 588532 268398 588768 268634
rect 588852 268398 589088 268634
rect 588532 232718 588768 232954
rect 588852 232718 589088 232954
rect 588532 232398 588768 232634
rect 588852 232398 589088 232634
rect 588532 196718 588768 196954
rect 588852 196718 589088 196954
rect 588532 196398 588768 196634
rect 588852 196398 589088 196634
rect 588532 160718 588768 160954
rect 588852 160718 589088 160954
rect 588532 160398 588768 160634
rect 588852 160398 589088 160634
rect 588532 124718 588768 124954
rect 588852 124718 589088 124954
rect 588532 124398 588768 124634
rect 588852 124398 589088 124634
rect 588532 88718 588768 88954
rect 588852 88718 589088 88954
rect 588532 88398 588768 88634
rect 588852 88398 589088 88634
rect 588532 52718 588768 52954
rect 588852 52718 589088 52954
rect 588532 52398 588768 52634
rect 588852 52398 589088 52634
rect 588532 16718 588768 16954
rect 588852 16718 589088 16954
rect 588532 16398 588768 16634
rect 588852 16398 589088 16634
rect 588532 -3772 588768 -3536
rect 588852 -3772 589088 -3536
rect 588532 -4092 588768 -3856
rect 588852 -4092 589088 -3856
rect 589492 669218 589728 669454
rect 589812 669218 590048 669454
rect 589492 668898 589728 669134
rect 589812 668898 590048 669134
rect 589492 633218 589728 633454
rect 589812 633218 590048 633454
rect 589492 632898 589728 633134
rect 589812 632898 590048 633134
rect 589492 597218 589728 597454
rect 589812 597218 590048 597454
rect 589492 596898 589728 597134
rect 589812 596898 590048 597134
rect 589492 561218 589728 561454
rect 589812 561218 590048 561454
rect 589492 560898 589728 561134
rect 589812 560898 590048 561134
rect 589492 525218 589728 525454
rect 589812 525218 590048 525454
rect 589492 524898 589728 525134
rect 589812 524898 590048 525134
rect 589492 489218 589728 489454
rect 589812 489218 590048 489454
rect 589492 488898 589728 489134
rect 589812 488898 590048 489134
rect 589492 453218 589728 453454
rect 589812 453218 590048 453454
rect 589492 452898 589728 453134
rect 589812 452898 590048 453134
rect 589492 417218 589728 417454
rect 589812 417218 590048 417454
rect 589492 416898 589728 417134
rect 589812 416898 590048 417134
rect 589492 381218 589728 381454
rect 589812 381218 590048 381454
rect 589492 380898 589728 381134
rect 589812 380898 590048 381134
rect 589492 345218 589728 345454
rect 589812 345218 590048 345454
rect 589492 344898 589728 345134
rect 589812 344898 590048 345134
rect 589492 309218 589728 309454
rect 589812 309218 590048 309454
rect 589492 308898 589728 309134
rect 589812 308898 590048 309134
rect 589492 273218 589728 273454
rect 589812 273218 590048 273454
rect 589492 272898 589728 273134
rect 589812 272898 590048 273134
rect 589492 237218 589728 237454
rect 589812 237218 590048 237454
rect 589492 236898 589728 237134
rect 589812 236898 590048 237134
rect 589492 201218 589728 201454
rect 589812 201218 590048 201454
rect 589492 200898 589728 201134
rect 589812 200898 590048 201134
rect 589492 165218 589728 165454
rect 589812 165218 590048 165454
rect 589492 164898 589728 165134
rect 589812 164898 590048 165134
rect 589492 129218 589728 129454
rect 589812 129218 590048 129454
rect 589492 128898 589728 129134
rect 589812 128898 590048 129134
rect 589492 93218 589728 93454
rect 589812 93218 590048 93454
rect 589492 92898 589728 93134
rect 589812 92898 590048 93134
rect 589492 57218 589728 57454
rect 589812 57218 590048 57454
rect 589492 56898 589728 57134
rect 589812 56898 590048 57134
rect 589492 21218 589728 21454
rect 589812 21218 590048 21454
rect 589492 20898 589728 21134
rect 589812 20898 590048 21134
rect 589492 -4732 589728 -4496
rect 589812 -4732 590048 -4496
rect 589492 -5052 589728 -4816
rect 589812 -5052 590048 -4816
rect 590452 673718 590688 673954
rect 590772 673718 591008 673954
rect 590452 673398 590688 673634
rect 590772 673398 591008 673634
rect 590452 637718 590688 637954
rect 590772 637718 591008 637954
rect 590452 637398 590688 637634
rect 590772 637398 591008 637634
rect 590452 601718 590688 601954
rect 590772 601718 591008 601954
rect 590452 601398 590688 601634
rect 590772 601398 591008 601634
rect 590452 565718 590688 565954
rect 590772 565718 591008 565954
rect 590452 565398 590688 565634
rect 590772 565398 591008 565634
rect 590452 529718 590688 529954
rect 590772 529718 591008 529954
rect 590452 529398 590688 529634
rect 590772 529398 591008 529634
rect 590452 493718 590688 493954
rect 590772 493718 591008 493954
rect 590452 493398 590688 493634
rect 590772 493398 591008 493634
rect 590452 457718 590688 457954
rect 590772 457718 591008 457954
rect 590452 457398 590688 457634
rect 590772 457398 591008 457634
rect 590452 421718 590688 421954
rect 590772 421718 591008 421954
rect 590452 421398 590688 421634
rect 590772 421398 591008 421634
rect 590452 385718 590688 385954
rect 590772 385718 591008 385954
rect 590452 385398 590688 385634
rect 590772 385398 591008 385634
rect 590452 349718 590688 349954
rect 590772 349718 591008 349954
rect 590452 349398 590688 349634
rect 590772 349398 591008 349634
rect 590452 313718 590688 313954
rect 590772 313718 591008 313954
rect 590452 313398 590688 313634
rect 590772 313398 591008 313634
rect 590452 277718 590688 277954
rect 590772 277718 591008 277954
rect 590452 277398 590688 277634
rect 590772 277398 591008 277634
rect 590452 241718 590688 241954
rect 590772 241718 591008 241954
rect 590452 241398 590688 241634
rect 590772 241398 591008 241634
rect 590452 205718 590688 205954
rect 590772 205718 591008 205954
rect 590452 205398 590688 205634
rect 590772 205398 591008 205634
rect 590452 169718 590688 169954
rect 590772 169718 591008 169954
rect 590452 169398 590688 169634
rect 590772 169398 591008 169634
rect 590452 133718 590688 133954
rect 590772 133718 591008 133954
rect 590452 133398 590688 133634
rect 590772 133398 591008 133634
rect 590452 97718 590688 97954
rect 590772 97718 591008 97954
rect 590452 97398 590688 97634
rect 590772 97398 591008 97634
rect 590452 61718 590688 61954
rect 590772 61718 591008 61954
rect 590452 61398 590688 61634
rect 590772 61398 591008 61634
rect 590452 25718 590688 25954
rect 590772 25718 591008 25954
rect 590452 25398 590688 25634
rect 590772 25398 591008 25634
rect 590452 -5692 590688 -5456
rect 590772 -5692 591008 -5456
rect 590452 -6012 590688 -5776
rect 590772 -6012 591008 -5776
rect 591412 678218 591648 678454
rect 591732 678218 591968 678454
rect 591412 677898 591648 678134
rect 591732 677898 591968 678134
rect 591412 642218 591648 642454
rect 591732 642218 591968 642454
rect 591412 641898 591648 642134
rect 591732 641898 591968 642134
rect 591412 606218 591648 606454
rect 591732 606218 591968 606454
rect 591412 605898 591648 606134
rect 591732 605898 591968 606134
rect 591412 570218 591648 570454
rect 591732 570218 591968 570454
rect 591412 569898 591648 570134
rect 591732 569898 591968 570134
rect 591412 534218 591648 534454
rect 591732 534218 591968 534454
rect 591412 533898 591648 534134
rect 591732 533898 591968 534134
rect 591412 498218 591648 498454
rect 591732 498218 591968 498454
rect 591412 497898 591648 498134
rect 591732 497898 591968 498134
rect 591412 462218 591648 462454
rect 591732 462218 591968 462454
rect 591412 461898 591648 462134
rect 591732 461898 591968 462134
rect 591412 426218 591648 426454
rect 591732 426218 591968 426454
rect 591412 425898 591648 426134
rect 591732 425898 591968 426134
rect 591412 390218 591648 390454
rect 591732 390218 591968 390454
rect 591412 389898 591648 390134
rect 591732 389898 591968 390134
rect 591412 354218 591648 354454
rect 591732 354218 591968 354454
rect 591412 353898 591648 354134
rect 591732 353898 591968 354134
rect 591412 318218 591648 318454
rect 591732 318218 591968 318454
rect 591412 317898 591648 318134
rect 591732 317898 591968 318134
rect 591412 282218 591648 282454
rect 591732 282218 591968 282454
rect 591412 281898 591648 282134
rect 591732 281898 591968 282134
rect 591412 246218 591648 246454
rect 591732 246218 591968 246454
rect 591412 245898 591648 246134
rect 591732 245898 591968 246134
rect 591412 210218 591648 210454
rect 591732 210218 591968 210454
rect 591412 209898 591648 210134
rect 591732 209898 591968 210134
rect 591412 174218 591648 174454
rect 591732 174218 591968 174454
rect 591412 173898 591648 174134
rect 591732 173898 591968 174134
rect 591412 138218 591648 138454
rect 591732 138218 591968 138454
rect 591412 137898 591648 138134
rect 591732 137898 591968 138134
rect 591412 102218 591648 102454
rect 591732 102218 591968 102454
rect 591412 101898 591648 102134
rect 591732 101898 591968 102134
rect 591412 66218 591648 66454
rect 591732 66218 591968 66454
rect 591412 65898 591648 66134
rect 591732 65898 591968 66134
rect 591412 30218 591648 30454
rect 591732 30218 591968 30454
rect 591412 29898 591648 30134
rect 591732 29898 591968 30134
rect 591412 -6652 591648 -6416
rect 591732 -6652 591968 -6416
rect 591412 -6972 591648 -6736
rect 591732 -6972 591968 -6736
rect 592372 682718 592608 682954
rect 592692 682718 592928 682954
rect 592372 682398 592608 682634
rect 592692 682398 592928 682634
rect 592372 646718 592608 646954
rect 592692 646718 592928 646954
rect 592372 646398 592608 646634
rect 592692 646398 592928 646634
rect 592372 610718 592608 610954
rect 592692 610718 592928 610954
rect 592372 610398 592608 610634
rect 592692 610398 592928 610634
rect 592372 574718 592608 574954
rect 592692 574718 592928 574954
rect 592372 574398 592608 574634
rect 592692 574398 592928 574634
rect 592372 538718 592608 538954
rect 592692 538718 592928 538954
rect 592372 538398 592608 538634
rect 592692 538398 592928 538634
rect 592372 502718 592608 502954
rect 592692 502718 592928 502954
rect 592372 502398 592608 502634
rect 592692 502398 592928 502634
rect 592372 466718 592608 466954
rect 592692 466718 592928 466954
rect 592372 466398 592608 466634
rect 592692 466398 592928 466634
rect 592372 430718 592608 430954
rect 592692 430718 592928 430954
rect 592372 430398 592608 430634
rect 592692 430398 592928 430634
rect 592372 394718 592608 394954
rect 592692 394718 592928 394954
rect 592372 394398 592608 394634
rect 592692 394398 592928 394634
rect 592372 358718 592608 358954
rect 592692 358718 592928 358954
rect 592372 358398 592608 358634
rect 592692 358398 592928 358634
rect 592372 322718 592608 322954
rect 592692 322718 592928 322954
rect 592372 322398 592608 322634
rect 592692 322398 592928 322634
rect 592372 286718 592608 286954
rect 592692 286718 592928 286954
rect 592372 286398 592608 286634
rect 592692 286398 592928 286634
rect 592372 250718 592608 250954
rect 592692 250718 592928 250954
rect 592372 250398 592608 250634
rect 592692 250398 592928 250634
rect 592372 214718 592608 214954
rect 592692 214718 592928 214954
rect 592372 214398 592608 214634
rect 592692 214398 592928 214634
rect 592372 178718 592608 178954
rect 592692 178718 592928 178954
rect 592372 178398 592608 178634
rect 592692 178398 592928 178634
rect 592372 142718 592608 142954
rect 592692 142718 592928 142954
rect 592372 142398 592608 142634
rect 592692 142398 592928 142634
rect 592372 106718 592608 106954
rect 592692 106718 592928 106954
rect 592372 106398 592608 106634
rect 592692 106398 592928 106634
rect 592372 70718 592608 70954
rect 592692 70718 592928 70954
rect 592372 70398 592608 70634
rect 592692 70398 592928 70634
rect 592372 34718 592608 34954
rect 592692 34718 592928 34954
rect 592372 34398 592608 34634
rect 592692 34398 592928 34634
rect 592372 -7612 592608 -7376
rect 592692 -7612 592928 -7376
rect 592372 -7932 592608 -7696
rect 592692 -7932 592928 -7696
<< metal5 >>
rect -9036 711868 592960 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect -9036 711548 592960 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect -9036 711280 592960 711312
rect -8076 710908 592000 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect -8076 710588 592000 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect -8076 710320 592000 710352
rect -7116 709948 591040 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect -7116 709628 591040 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect -7116 709360 591040 709392
rect -6156 708988 590080 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect -6156 708668 590080 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect -6156 708400 590080 708432
rect -5196 708028 589120 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect -5196 707708 589120 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect -5196 707440 589120 707472
rect -4236 707068 588160 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect -4236 706748 588160 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect -4236 706480 588160 706512
rect -3276 706108 587200 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect -3276 705788 587200 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect -3276 705520 587200 705552
rect -2316 705148 586240 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect -2316 704828 586240 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect -2316 704560 586240 704592
rect -9036 700954 592960 700986
rect -9036 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 592960 700954
rect -9036 700634 592960 700718
rect -9036 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 592960 700634
rect -9036 700366 592960 700398
rect -9036 696454 592960 696486
rect -9036 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 592960 696454
rect -9036 696134 592960 696218
rect -9036 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 592960 696134
rect -9036 695866 592960 695898
rect -9036 691954 592960 691986
rect -9036 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 592960 691954
rect -9036 691634 592960 691718
rect -9036 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 592960 691634
rect -9036 691366 592960 691398
rect -9036 687454 592960 687486
rect -9036 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 592960 687454
rect -9036 687134 592960 687218
rect -9036 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 592960 687134
rect -9036 686866 592960 686898
rect -9036 682954 592960 682986
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect -9036 682634 592960 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect -9036 682366 592960 682398
rect -9036 678454 592960 678486
rect -9036 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592960 678454
rect -9036 678134 592960 678218
rect -9036 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592960 678134
rect -9036 677866 592960 677898
rect -9036 673954 592960 673986
rect -9036 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 592960 673954
rect -9036 673634 592960 673718
rect -9036 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 592960 673634
rect -9036 673366 592960 673398
rect -9036 669454 592960 669486
rect -9036 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 592960 669454
rect -9036 669134 592960 669218
rect -9036 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 592960 669134
rect -9036 668866 592960 668898
rect -9036 664954 592960 664986
rect -9036 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 592960 664954
rect -9036 664634 592960 664718
rect -9036 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 592960 664634
rect -9036 664366 592960 664398
rect -9036 660454 592960 660486
rect -9036 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 592960 660454
rect -9036 660134 592960 660218
rect -9036 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 592960 660134
rect -9036 659866 592960 659898
rect -9036 655954 592960 655986
rect -9036 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 592960 655954
rect -9036 655634 592960 655718
rect -9036 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 592960 655634
rect -9036 655366 592960 655398
rect -9036 651454 592960 651486
rect -9036 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 592960 651454
rect -9036 651134 592960 651218
rect -9036 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 592960 651134
rect -9036 650866 592960 650898
rect -9036 646954 592960 646986
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect -9036 646634 592960 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect -9036 646366 592960 646398
rect -9036 642454 592960 642486
rect -9036 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592960 642454
rect -9036 642134 592960 642218
rect -9036 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592960 642134
rect -9036 641866 592960 641898
rect -9036 637954 592960 637986
rect -9036 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 592960 637954
rect -9036 637634 592960 637718
rect -9036 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 592960 637634
rect -9036 637366 592960 637398
rect -9036 633454 592960 633486
rect -9036 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 592960 633454
rect -9036 633134 592960 633218
rect -9036 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 592960 633134
rect -9036 632866 592960 632898
rect -9036 628954 592960 628986
rect -9036 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 592960 628954
rect -9036 628634 592960 628718
rect -9036 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 592960 628634
rect -9036 628366 592960 628398
rect -9036 624454 592960 624486
rect -9036 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 592960 624454
rect -9036 624134 592960 624218
rect -9036 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 592960 624134
rect -9036 623866 592960 623898
rect -9036 619954 592960 619986
rect -9036 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 592960 619954
rect -9036 619634 592960 619718
rect -9036 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 592960 619634
rect -9036 619366 592960 619398
rect -9036 615454 592960 615486
rect -9036 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 592960 615454
rect -9036 615134 592960 615218
rect -9036 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 592960 615134
rect -9036 614866 592960 614898
rect -9036 610954 592960 610986
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect -9036 610634 592960 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect -9036 610366 592960 610398
rect -9036 606454 592960 606486
rect -9036 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592960 606454
rect -9036 606134 592960 606218
rect -9036 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592960 606134
rect -9036 605866 592960 605898
rect -9036 601954 592960 601986
rect -9036 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 592960 601954
rect -9036 601634 592960 601718
rect -9036 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 592960 601634
rect -9036 601366 592960 601398
rect -9036 597454 592960 597486
rect -9036 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 592960 597454
rect -9036 597134 592960 597218
rect -9036 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 592960 597134
rect -9036 596866 592960 596898
rect -9036 592954 592960 592986
rect -9036 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 592960 592954
rect -9036 592634 592960 592718
rect -9036 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 592960 592634
rect -9036 592366 592960 592398
rect -9036 588454 592960 588486
rect -9036 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 592960 588454
rect -9036 588134 592960 588218
rect -9036 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 592960 588134
rect -9036 587866 592960 587898
rect -9036 583954 592960 583986
rect -9036 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 592960 583954
rect -9036 583634 592960 583718
rect -9036 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 592960 583634
rect -9036 583366 592960 583398
rect -9036 579454 592960 579486
rect -9036 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 592960 579454
rect -9036 579134 592960 579218
rect -9036 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 592960 579134
rect -9036 578866 592960 578898
rect -9036 574954 592960 574986
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect -9036 574634 592960 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect -9036 574366 592960 574398
rect -9036 570454 592960 570486
rect -9036 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592960 570454
rect -9036 570134 592960 570218
rect -9036 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592960 570134
rect -9036 569866 592960 569898
rect -9036 565954 592960 565986
rect -9036 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 592960 565954
rect -9036 565634 592960 565718
rect -9036 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 592960 565634
rect -9036 565366 592960 565398
rect -9036 561454 592960 561486
rect -9036 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 592960 561454
rect -9036 561134 592960 561218
rect -9036 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 592960 561134
rect -9036 560866 592960 560898
rect -9036 556954 592960 556986
rect -9036 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 592960 556954
rect -9036 556634 592960 556718
rect -9036 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 592960 556634
rect -9036 556366 592960 556398
rect -9036 552454 592960 552486
rect -9036 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 592960 552454
rect -9036 552134 592960 552218
rect -9036 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 592960 552134
rect -9036 551866 592960 551898
rect -9036 547954 592960 547986
rect -9036 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 592960 547954
rect -9036 547634 592960 547718
rect -9036 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 592960 547634
rect -9036 547366 592960 547398
rect -9036 543454 592960 543486
rect -9036 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 592960 543454
rect -9036 543134 592960 543218
rect -9036 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 592960 543134
rect -9036 542866 592960 542898
rect -9036 538954 592960 538986
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect -9036 538634 592960 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect -9036 538366 592960 538398
rect -9036 534454 592960 534486
rect -9036 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592960 534454
rect -9036 534134 592960 534218
rect -9036 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592960 534134
rect -9036 533866 592960 533898
rect -9036 529954 592960 529986
rect -9036 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 592960 529954
rect -9036 529634 592960 529718
rect -9036 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 592960 529634
rect -9036 529366 592960 529398
rect -9036 525454 592960 525486
rect -9036 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 592960 525454
rect -9036 525134 592960 525218
rect -9036 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 592960 525134
rect -9036 524866 592960 524898
rect -9036 520954 592960 520986
rect -9036 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 592960 520954
rect -9036 520634 592960 520718
rect -9036 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 592960 520634
rect -9036 520366 592960 520398
rect -9036 516454 592960 516486
rect -9036 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 592960 516454
rect -9036 516134 592960 516218
rect -9036 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 592960 516134
rect -9036 515866 592960 515898
rect -9036 511954 592960 511986
rect -9036 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 592960 511954
rect -9036 511634 592960 511718
rect -9036 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 592960 511634
rect -9036 511366 592960 511398
rect -9036 507454 592960 507486
rect -9036 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 592960 507454
rect -9036 507134 592960 507218
rect -9036 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 592960 507134
rect -9036 506866 592960 506898
rect -9036 502954 592960 502986
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect -9036 502634 592960 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect -9036 502366 592960 502398
rect -9036 498454 592960 498486
rect -9036 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592960 498454
rect -9036 498134 592960 498218
rect -9036 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592960 498134
rect -9036 497866 592960 497898
rect -9036 493954 592960 493986
rect -9036 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 592960 493954
rect -9036 493634 592960 493718
rect -9036 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 592960 493634
rect -9036 493366 592960 493398
rect -9036 489454 592960 489486
rect -9036 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 592960 489454
rect -9036 489134 592960 489218
rect -9036 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 592960 489134
rect -9036 488866 592960 488898
rect -9036 484954 592960 484986
rect -9036 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 592960 484954
rect -9036 484634 592960 484718
rect -9036 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 592960 484634
rect -9036 484366 592960 484398
rect -9036 480454 592960 480486
rect -9036 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 592960 480454
rect -9036 480134 592960 480218
rect -9036 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 592960 480134
rect -9036 479866 592960 479898
rect -9036 475954 592960 475986
rect -9036 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 592960 475954
rect -9036 475634 592960 475718
rect -9036 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 592960 475634
rect -9036 475366 592960 475398
rect -9036 471454 592960 471486
rect -9036 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 592960 471454
rect -9036 471134 592960 471218
rect -9036 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 592960 471134
rect -9036 470866 592960 470898
rect -9036 466954 592960 466986
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect -9036 466634 592960 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect -9036 466366 592960 466398
rect -9036 462454 592960 462486
rect -9036 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592960 462454
rect -9036 462134 592960 462218
rect -9036 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592960 462134
rect -9036 461866 592960 461898
rect -9036 457954 592960 457986
rect -9036 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 592960 457954
rect -9036 457634 592960 457718
rect -9036 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 592960 457634
rect -9036 457366 592960 457398
rect -9036 453454 592960 453486
rect -9036 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 592960 453454
rect -9036 453134 592960 453218
rect -9036 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 592960 453134
rect -9036 452866 592960 452898
rect -9036 448954 592960 448986
rect -9036 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 592960 448954
rect -9036 448634 592960 448718
rect -9036 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 592960 448634
rect -9036 448366 592960 448398
rect -9036 444454 592960 444486
rect -9036 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 592960 444454
rect -9036 444134 592960 444218
rect -9036 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 592960 444134
rect -9036 443866 592960 443898
rect -9036 439954 592960 439986
rect -9036 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 592960 439954
rect -9036 439634 592960 439718
rect -9036 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 592960 439634
rect -9036 439366 592960 439398
rect -9036 435454 592960 435486
rect -9036 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 592960 435454
rect -9036 435134 592960 435218
rect -9036 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 592960 435134
rect -9036 434866 592960 434898
rect -9036 430954 592960 430986
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect -9036 430634 592960 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect -9036 430366 592960 430398
rect -9036 426454 592960 426486
rect -9036 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592960 426454
rect -9036 426134 592960 426218
rect -9036 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592960 426134
rect -9036 425866 592960 425898
rect -9036 421954 592960 421986
rect -9036 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 592960 421954
rect -9036 421634 592960 421718
rect -9036 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 592960 421634
rect -9036 421366 592960 421398
rect -9036 417454 592960 417486
rect -9036 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 592960 417454
rect -9036 417134 592960 417218
rect -9036 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 592960 417134
rect -9036 416866 592960 416898
rect -9036 412954 592960 412986
rect -9036 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 592960 412954
rect -9036 412634 592960 412718
rect -9036 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 592960 412634
rect -9036 412366 592960 412398
rect -9036 408454 592960 408486
rect -9036 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 592960 408454
rect -9036 408134 592960 408218
rect -9036 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 592960 408134
rect -9036 407866 592960 407898
rect -9036 403954 592960 403986
rect -9036 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 592960 403954
rect -9036 403634 592960 403718
rect -9036 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 592960 403634
rect -9036 403366 592960 403398
rect -9036 399454 592960 399486
rect -9036 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 592960 399454
rect -9036 399134 592960 399218
rect -9036 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 592960 399134
rect -9036 398866 592960 398898
rect -9036 394954 592960 394986
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect -9036 394634 592960 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect -9036 394366 592960 394398
rect -9036 390454 592960 390486
rect -9036 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592960 390454
rect -9036 390134 592960 390218
rect -9036 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592960 390134
rect -9036 389866 592960 389898
rect -9036 385954 592960 385986
rect -9036 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 592960 385954
rect -9036 385634 592960 385718
rect -9036 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 592960 385634
rect -9036 385366 592960 385398
rect -9036 381454 592960 381486
rect -9036 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 592960 381454
rect -9036 381134 592960 381218
rect -9036 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 592960 381134
rect -9036 380866 592960 380898
rect -9036 376954 592960 376986
rect -9036 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 592960 376954
rect -9036 376634 592960 376718
rect -9036 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 592960 376634
rect -9036 376366 592960 376398
rect -9036 372454 592960 372486
rect -9036 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 592960 372454
rect -9036 372134 592960 372218
rect -9036 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 592960 372134
rect -9036 371866 592960 371898
rect -9036 367954 592960 367986
rect -9036 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 592960 367954
rect -9036 367634 592960 367718
rect -9036 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 592960 367634
rect -9036 367366 592960 367398
rect -9036 363454 592960 363486
rect -9036 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 592960 363454
rect -9036 363134 592960 363218
rect -9036 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 592960 363134
rect -9036 362866 592960 362898
rect -9036 358954 592960 358986
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect -9036 358634 592960 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect -9036 358366 592960 358398
rect -9036 354454 592960 354486
rect -9036 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592960 354454
rect -9036 354134 592960 354218
rect -9036 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592960 354134
rect -9036 353866 592960 353898
rect -9036 349954 592960 349986
rect -9036 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 592960 349954
rect -9036 349634 592960 349718
rect -9036 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 592960 349634
rect -9036 349366 592960 349398
rect -9036 345454 592960 345486
rect -9036 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 592960 345454
rect -9036 345134 592960 345218
rect -9036 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 592960 345134
rect -9036 344866 592960 344898
rect -9036 340954 592960 340986
rect -9036 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 592960 340954
rect -9036 340634 592960 340718
rect -9036 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 592960 340634
rect -9036 340366 592960 340398
rect -9036 336454 592960 336486
rect -9036 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 592960 336454
rect -9036 336134 592960 336218
rect -9036 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 592960 336134
rect -9036 335866 592960 335898
rect -9036 331954 592960 331986
rect -9036 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 592960 331954
rect -9036 331634 592960 331718
rect -9036 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 592960 331634
rect -9036 331366 592960 331398
rect -9036 327454 592960 327486
rect -9036 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 592960 327454
rect -9036 327134 592960 327218
rect -9036 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 592960 327134
rect -9036 326866 592960 326898
rect -9036 322954 592960 322986
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect -9036 322634 592960 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect -9036 322366 592960 322398
rect -9036 318454 592960 318486
rect -9036 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592960 318454
rect -9036 318134 592960 318218
rect -9036 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592960 318134
rect -9036 317866 592960 317898
rect -9036 313954 592960 313986
rect -9036 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 592960 313954
rect -9036 313634 592960 313718
rect -9036 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 592960 313634
rect -9036 313366 592960 313398
rect -9036 309454 592960 309486
rect -9036 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 592960 309454
rect -9036 309134 592960 309218
rect -9036 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 592960 309134
rect -9036 308866 592960 308898
rect -9036 304954 592960 304986
rect -9036 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 592960 304954
rect -9036 304634 592960 304718
rect -9036 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 592960 304634
rect -9036 304366 592960 304398
rect -9036 300454 592960 300486
rect -9036 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 592960 300454
rect -9036 300134 592960 300218
rect -9036 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 592960 300134
rect -9036 299866 592960 299898
rect -9036 295954 592960 295986
rect -9036 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 592960 295954
rect -9036 295634 592960 295718
rect -9036 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 592960 295634
rect -9036 295366 592960 295398
rect -9036 291454 592960 291486
rect -9036 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 592960 291454
rect -9036 291134 592960 291218
rect -9036 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 592960 291134
rect -9036 290866 592960 290898
rect -9036 286954 592960 286986
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect -9036 286634 592960 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect -9036 286366 592960 286398
rect -9036 282454 592960 282486
rect -9036 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592960 282454
rect -9036 282134 592960 282218
rect -9036 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592960 282134
rect -9036 281866 592960 281898
rect -9036 277954 592960 277986
rect -9036 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 592960 277954
rect -9036 277634 592960 277718
rect -9036 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 592960 277634
rect -9036 277366 592960 277398
rect -9036 273454 592960 273486
rect -9036 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 592960 273454
rect -9036 273134 592960 273218
rect -9036 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 592960 273134
rect -9036 272866 592960 272898
rect -9036 268954 592960 268986
rect -9036 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 592960 268954
rect -9036 268634 592960 268718
rect -9036 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 592960 268634
rect -9036 268366 592960 268398
rect -9036 264454 592960 264486
rect -9036 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 592960 264454
rect -9036 264134 592960 264218
rect -9036 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 592960 264134
rect -9036 263866 592960 263898
rect -9036 259954 592960 259986
rect -9036 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 592960 259954
rect -9036 259634 592960 259718
rect -9036 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 592960 259634
rect -9036 259366 592960 259398
rect -9036 255454 592960 255486
rect -9036 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 236250 255454
rect 236486 255218 266970 255454
rect 267206 255218 297690 255454
rect 297926 255218 328410 255454
rect 328646 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 592960 255454
rect -9036 255134 592960 255218
rect -9036 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 236250 255134
rect 236486 254898 266970 255134
rect 267206 254898 297690 255134
rect 297926 254898 328410 255134
rect 328646 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 592960 255134
rect -9036 254866 592960 254898
rect -9036 250954 592960 250986
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect -9036 250634 592960 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect -9036 250366 592960 250398
rect -9036 246454 592960 246486
rect -9036 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592960 246454
rect -9036 246134 592960 246218
rect -9036 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592960 246134
rect -9036 245866 592960 245898
rect -9036 241954 592960 241986
rect -9036 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 592960 241954
rect -9036 241634 592960 241718
rect -9036 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 592960 241634
rect -9036 241366 592960 241398
rect -9036 237454 592960 237486
rect -9036 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 592960 237454
rect -9036 237134 592960 237218
rect -9036 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 592960 237134
rect -9036 236866 592960 236898
rect -9036 232954 592960 232986
rect -9036 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 592960 232954
rect -9036 232634 592960 232718
rect -9036 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 592960 232634
rect -9036 232366 592960 232398
rect -9036 228454 592960 228486
rect -9036 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 592960 228454
rect -9036 228134 592960 228218
rect -9036 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 592960 228134
rect -9036 227866 592960 227898
rect -9036 223954 592960 223986
rect -9036 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 251610 223954
rect 251846 223718 282330 223954
rect 282566 223718 313050 223954
rect 313286 223718 343770 223954
rect 344006 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 592960 223954
rect -9036 223634 592960 223718
rect -9036 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 251610 223634
rect 251846 223398 282330 223634
rect 282566 223398 313050 223634
rect 313286 223398 343770 223634
rect 344006 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 592960 223634
rect -9036 223366 592960 223398
rect -9036 219454 592960 219486
rect -9036 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 236250 219454
rect 236486 219218 266970 219454
rect 267206 219218 297690 219454
rect 297926 219218 328410 219454
rect 328646 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 592960 219454
rect -9036 219134 592960 219218
rect -9036 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 236250 219134
rect 236486 218898 266970 219134
rect 267206 218898 297690 219134
rect 297926 218898 328410 219134
rect 328646 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 592960 219134
rect -9036 218866 592960 218898
rect -9036 214954 592960 214986
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect -9036 214634 592960 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect -9036 214366 592960 214398
rect -9036 210454 592960 210486
rect -9036 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592960 210454
rect -9036 210134 592960 210218
rect -9036 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592960 210134
rect -9036 209866 592960 209898
rect -9036 205954 592960 205986
rect -9036 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 592960 205954
rect -9036 205634 592960 205718
rect -9036 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 592960 205634
rect -9036 205366 592960 205398
rect -9036 201454 592960 201486
rect -9036 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 592960 201454
rect -9036 201134 592960 201218
rect -9036 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 592960 201134
rect -9036 200866 592960 200898
rect -9036 196954 592960 196986
rect -9036 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 592960 196954
rect -9036 196634 592960 196718
rect -9036 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 592960 196634
rect -9036 196366 592960 196398
rect -9036 192454 592960 192486
rect -9036 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 592960 192454
rect -9036 192134 592960 192218
rect -9036 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 592960 192134
rect -9036 191866 592960 191898
rect -9036 187954 592960 187986
rect -9036 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 251610 187954
rect 251846 187718 282330 187954
rect 282566 187718 313050 187954
rect 313286 187718 343770 187954
rect 344006 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 592960 187954
rect -9036 187634 592960 187718
rect -9036 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 251610 187634
rect 251846 187398 282330 187634
rect 282566 187398 313050 187634
rect 313286 187398 343770 187634
rect 344006 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 592960 187634
rect -9036 187366 592960 187398
rect -9036 183454 592960 183486
rect -9036 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 236250 183454
rect 236486 183218 266970 183454
rect 267206 183218 297690 183454
rect 297926 183218 328410 183454
rect 328646 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 592960 183454
rect -9036 183134 592960 183218
rect -9036 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 236250 183134
rect 236486 182898 266970 183134
rect 267206 182898 297690 183134
rect 297926 182898 328410 183134
rect 328646 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 592960 183134
rect -9036 182866 592960 182898
rect -9036 178954 592960 178986
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect -9036 178634 592960 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect -9036 178366 592960 178398
rect -9036 174454 592960 174486
rect -9036 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592960 174454
rect -9036 174134 592960 174218
rect -9036 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592960 174134
rect -9036 173866 592960 173898
rect -9036 169954 592960 169986
rect -9036 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 592960 169954
rect -9036 169634 592960 169718
rect -9036 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 592960 169634
rect -9036 169366 592960 169398
rect -9036 165454 592960 165486
rect -9036 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 592960 165454
rect -9036 165134 592960 165218
rect -9036 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 592960 165134
rect -9036 164866 592960 164898
rect -9036 160954 592960 160986
rect -9036 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 592960 160954
rect -9036 160634 592960 160718
rect -9036 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 592960 160634
rect -9036 160366 592960 160398
rect -9036 156454 592960 156486
rect -9036 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 592960 156454
rect -9036 156134 592960 156218
rect -9036 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 592960 156134
rect -9036 155866 592960 155898
rect -9036 151954 592960 151986
rect -9036 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 251610 151954
rect 251846 151718 282330 151954
rect 282566 151718 313050 151954
rect 313286 151718 343770 151954
rect 344006 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 592960 151954
rect -9036 151634 592960 151718
rect -9036 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 251610 151634
rect 251846 151398 282330 151634
rect 282566 151398 313050 151634
rect 313286 151398 343770 151634
rect 344006 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 592960 151634
rect -9036 151366 592960 151398
rect -9036 147454 592960 147486
rect -9036 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 236250 147454
rect 236486 147218 266970 147454
rect 267206 147218 297690 147454
rect 297926 147218 328410 147454
rect 328646 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 592960 147454
rect -9036 147134 592960 147218
rect -9036 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 236250 147134
rect 236486 146898 266970 147134
rect 267206 146898 297690 147134
rect 297926 146898 328410 147134
rect 328646 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 592960 147134
rect -9036 146866 592960 146898
rect -9036 142954 592960 142986
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect -9036 142634 592960 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect -9036 142366 592960 142398
rect -9036 138454 592960 138486
rect -9036 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592960 138454
rect -9036 138134 592960 138218
rect -9036 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592960 138134
rect -9036 137866 592960 137898
rect -9036 133954 592960 133986
rect -9036 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 592960 133954
rect -9036 133634 592960 133718
rect -9036 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 592960 133634
rect -9036 133366 592960 133398
rect -9036 129454 592960 129486
rect -9036 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 592960 129454
rect -9036 129134 592960 129218
rect -9036 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 592960 129134
rect -9036 128866 592960 128898
rect -9036 124954 592960 124986
rect -9036 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 592960 124954
rect -9036 124634 592960 124718
rect -9036 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 592960 124634
rect -9036 124366 592960 124398
rect -9036 120454 592960 120486
rect -9036 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 592960 120454
rect -9036 120134 592960 120218
rect -9036 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 592960 120134
rect -9036 119866 592960 119898
rect -9036 115954 592960 115986
rect -9036 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 251610 115954
rect 251846 115718 282330 115954
rect 282566 115718 313050 115954
rect 313286 115718 343770 115954
rect 344006 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 592960 115954
rect -9036 115634 592960 115718
rect -9036 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 251610 115634
rect 251846 115398 282330 115634
rect 282566 115398 313050 115634
rect 313286 115398 343770 115634
rect 344006 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 592960 115634
rect -9036 115366 592960 115398
rect -9036 111454 592960 111486
rect -9036 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 236250 111454
rect 236486 111218 266970 111454
rect 267206 111218 297690 111454
rect 297926 111218 328410 111454
rect 328646 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 592960 111454
rect -9036 111134 592960 111218
rect -9036 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 236250 111134
rect 236486 110898 266970 111134
rect 267206 110898 297690 111134
rect 297926 110898 328410 111134
rect 328646 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 592960 111134
rect -9036 110866 592960 110898
rect -9036 106954 592960 106986
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect -9036 106634 592960 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect -9036 106366 592960 106398
rect -9036 102454 592960 102486
rect -9036 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592960 102454
rect -9036 102134 592960 102218
rect -9036 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592960 102134
rect -9036 101866 592960 101898
rect -9036 97954 592960 97986
rect -9036 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 592960 97954
rect -9036 97634 592960 97718
rect -9036 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 592960 97634
rect -9036 97366 592960 97398
rect -9036 93454 592960 93486
rect -9036 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 592960 93454
rect -9036 93134 592960 93218
rect -9036 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 592960 93134
rect -9036 92866 592960 92898
rect -9036 88954 592960 88986
rect -9036 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 592960 88954
rect -9036 88634 592960 88718
rect -9036 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 592960 88634
rect -9036 88366 592960 88398
rect -9036 84454 592960 84486
rect -9036 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 592960 84454
rect -9036 84134 592960 84218
rect -9036 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 592960 84134
rect -9036 83866 592960 83898
rect -9036 79954 592960 79986
rect -9036 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 592960 79954
rect -9036 79634 592960 79718
rect -9036 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 592960 79634
rect -9036 79366 592960 79398
rect -9036 75454 592960 75486
rect -9036 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 592960 75454
rect -9036 75134 592960 75218
rect -9036 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 592960 75134
rect -9036 74866 592960 74898
rect -9036 70954 592960 70986
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect -9036 70634 592960 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect -9036 70366 592960 70398
rect -9036 66454 592960 66486
rect -9036 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592960 66454
rect -9036 66134 592960 66218
rect -9036 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592960 66134
rect -9036 65866 592960 65898
rect -9036 61954 592960 61986
rect -9036 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 592960 61954
rect -9036 61634 592960 61718
rect -9036 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 592960 61634
rect -9036 61366 592960 61398
rect -9036 57454 592960 57486
rect -9036 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 592960 57454
rect -9036 57134 592960 57218
rect -9036 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 592960 57134
rect -9036 56866 592960 56898
rect -9036 52954 592960 52986
rect -9036 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 592960 52954
rect -9036 52634 592960 52718
rect -9036 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 592960 52634
rect -9036 52366 592960 52398
rect -9036 48454 592960 48486
rect -9036 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 592960 48454
rect -9036 48134 592960 48218
rect -9036 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 592960 48134
rect -9036 47866 592960 47898
rect -9036 43954 592960 43986
rect -9036 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 592960 43954
rect -9036 43634 592960 43718
rect -9036 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 592960 43634
rect -9036 43366 592960 43398
rect -9036 39454 592960 39486
rect -9036 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 592960 39454
rect -9036 39134 592960 39218
rect -9036 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 592960 39134
rect -9036 38866 592960 38898
rect -9036 34954 592960 34986
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect -9036 34634 592960 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect -9036 34366 592960 34398
rect -9036 30454 592960 30486
rect -9036 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592960 30454
rect -9036 30134 592960 30218
rect -9036 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592960 30134
rect -9036 29866 592960 29898
rect -9036 25954 592960 25986
rect -9036 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 592960 25954
rect -9036 25634 592960 25718
rect -9036 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 592960 25634
rect -9036 25366 592960 25398
rect -9036 21454 592960 21486
rect -9036 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 592960 21454
rect -9036 21134 592960 21218
rect -9036 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 592960 21134
rect -9036 20866 592960 20898
rect -9036 16954 592960 16986
rect -9036 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 592960 16954
rect -9036 16634 592960 16718
rect -9036 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 592960 16634
rect -9036 16366 592960 16398
rect -9036 12454 592960 12486
rect -9036 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 592960 12454
rect -9036 12134 592960 12218
rect -9036 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 592960 12134
rect -9036 11866 592960 11898
rect -9036 7954 592960 7986
rect -9036 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 592960 7954
rect -9036 7634 592960 7718
rect -9036 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 592960 7634
rect -9036 7366 592960 7398
rect -9036 3454 592960 3486
rect -9036 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 592960 3454
rect -9036 3134 592960 3218
rect -9036 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 592960 3134
rect -9036 2866 592960 2898
rect -2316 -656 586240 -624
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect -2316 -976 586240 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect -2316 -1244 586240 -1212
rect -3276 -1616 587200 -1584
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect -3276 -1936 587200 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect -3276 -2204 587200 -2172
rect -4236 -2576 588160 -2544
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect -4236 -2896 588160 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect -4236 -3164 588160 -3132
rect -5196 -3536 589120 -3504
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect -5196 -3856 589120 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect -5196 -4124 589120 -4092
rect -6156 -4496 590080 -4464
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect -6156 -4816 590080 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect -6156 -5084 590080 -5052
rect -7116 -5456 591040 -5424
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect -7116 -5776 591040 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect -7116 -6044 591040 -6012
rect -8076 -6416 592000 -6384
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect -8076 -6736 592000 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect -8076 -7004 592000 -6972
rect -9036 -7376 592960 -7344
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect -9036 -7696 592960 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect -9036 -7964 592960 -7932
use user_proj_example  mprj
timestamp 0
transform 1 0 232000 0 1 100000
box 0 0 120000 160000
<< labels >>
flabel metal3 s 583520 285820 584960 286060 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 445730 703520 445842 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 380962 703520 381074 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316194 703520 316306 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186658 703520 186770 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121890 703520 122002 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 57122 703520 57234 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 694228 480 694468 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 642548 480 642788 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 590868 480 591108 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338588 584960 338828 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 539188 480 539428 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 487508 480 487748 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 435828 480 436068 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384148 480 384388 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332468 480 332708 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 280788 480 281028 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 229108 480 229348 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 177428 480 177668 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 125748 480 125988 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391356 584960 391596 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444124 584960 444364 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 496892 584960 497132 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 549660 584960 549900 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 602428 584960 602668 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 655196 584960 655436 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575266 703520 575378 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510498 703520 510610 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 8788 584960 9028 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457316 584960 457556 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 510084 584960 510324 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 562852 584960 563092 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 615620 584960 615860 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 668388 584960 668628 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559074 703520 559186 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494306 703520 494418 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429538 703520 429650 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364770 703520 364882 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300002 703520 300114 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 48364 584960 48604 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235234 703520 235346 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170466 703520 170578 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105698 703520 105810 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40930 703520 41042 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 681308 480 681548 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 629628 480 629868 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 577948 480 578188 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 526268 480 526508 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 474588 480 474828 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 422908 480 423148 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 87940 584960 88180 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319548 480 319788 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267868 480 268108 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 216188 480 216428 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 164508 480 164748 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 112828 480 113068 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 74068 480 74308 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 35308 480 35548 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 127516 584960 127756 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 167092 584960 167332 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 206668 584960 206908 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 246244 584960 246484 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 299012 584960 299252 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404548 584960 404788 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 35172 584960 35412 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 483700 584960 483940 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 536468 584960 536708 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 589236 584960 589476 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 642004 584960 642244 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 694772 584960 695012 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 526690 703520 526802 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 461922 703520 462034 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397154 703520 397266 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332386 703520 332498 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 74748 584960 74988 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202850 703520 202962 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 138082 703520 138194 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 73314 703520 73426 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8546 703520 8658 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 655468 480 655708 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 603788 480 604028 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 552108 480 552348 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 500428 480 500668 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 448748 480 448988 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397068 480 397308 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 114324 584960 114564 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345388 480 345628 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293708 480 293948 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 242028 480 242268 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 190348 480 190588 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 138668 480 138908 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 86988 480 87228 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 48228 480 48468 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 9468 480 9708 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 153900 584960 154140 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 193476 584960 193716 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 233052 584960 233292 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272628 584960 272868 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325396 584960 325636 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378164 584960 378404 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 430932 584960 431172 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 21980 584960 22220 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 470508 584960 470748 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 523276 584960 523516 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 576044 584960 576284 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 628812 584960 629052 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 681580 584960 681820 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 542882 703520 542994 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478114 703520 478226 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413346 703520 413458 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348578 703520 348690 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 61556 584960 61796 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 219042 703520 219154 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154274 703520 154386 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89506 703520 89618 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24738 703520 24850 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 668388 480 668628 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 616708 480 616948 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 565028 480 565268 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 513348 480 513588 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 461668 480 461908 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 409988 480 410228 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 101132 584960 101372 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306628 480 306868 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 254948 480 255188 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 203268 480 203508 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 151588 480 151828 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 99908 480 100148 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 61148 480 61388 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 22388 480 22628 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 140708 584960 140948 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 180284 584960 180524 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 219860 584960 220100 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 259436 584960 259676 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 312204 584960 312444 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 417740 584960 417980 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 136794 -960 136906 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 467994 -960 468106 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 471306 -960 471418 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 474618 -960 474730 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 477930 -960 478042 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 481242 -960 481354 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 484554 -960 484666 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 487866 -960 487978 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 491178 -960 491290 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 494490 -960 494602 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 497802 -960 497914 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 169914 -960 170026 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 501114 -960 501226 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 504426 -960 504538 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 507738 -960 507850 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 511050 -960 511162 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 514362 -960 514474 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 517674 -960 517786 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 520986 -960 521098 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 524298 -960 524410 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 527610 -960 527722 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 530922 -960 531034 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 173226 -960 173338 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 534234 -960 534346 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 537546 -960 537658 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 540858 -960 540970 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 544170 -960 544282 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 547482 -960 547594 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 550794 -960 550906 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 554106 -960 554218 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 557418 -960 557530 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 176538 -960 176650 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 179850 -960 179962 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 183162 -960 183274 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 186474 -960 186586 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 189786 -960 189898 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 193098 -960 193210 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 196410 -960 196522 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 199722 -960 199834 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 140106 -960 140218 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 203034 -960 203146 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 206346 -960 206458 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 209658 -960 209770 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 212970 -960 213082 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 216282 -960 216394 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 219594 -960 219706 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 222906 -960 223018 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 226218 -960 226330 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 229530 -960 229642 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 232842 -960 232954 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 143418 -960 143530 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 236154 -960 236266 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 239466 -960 239578 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 242778 -960 242890 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 246090 -960 246202 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 249402 -960 249514 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 252714 -960 252826 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 256026 -960 256138 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 259338 -960 259450 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 262650 -960 262762 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 265962 -960 266074 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 146730 -960 146842 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 269274 -960 269386 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 272586 -960 272698 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 275898 -960 276010 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 279210 -960 279322 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 282522 -960 282634 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285834 -960 285946 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 289146 -960 289258 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292458 -960 292570 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 295770 -960 295882 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299082 -960 299194 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 150042 -960 150154 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 302394 -960 302506 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 305706 -960 305818 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 312330 -960 312442 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 315642 -960 315754 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 318954 -960 319066 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 322266 -960 322378 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 328890 -960 329002 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 332202 -960 332314 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 153354 -960 153466 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 335514 -960 335626 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 338826 -960 338938 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 345450 -960 345562 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 348762 -960 348874 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 352074 -960 352186 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 355386 -960 355498 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 362010 -960 362122 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 365322 -960 365434 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 156666 -960 156778 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 368634 -960 368746 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 371946 -960 372058 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 378570 -960 378682 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 381882 -960 381994 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 385194 -960 385306 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 388506 -960 388618 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 395130 -960 395242 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 398442 -960 398554 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 159978 -960 160090 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 401754 -960 401866 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 405066 -960 405178 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 411690 -960 411802 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 415002 -960 415114 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 418314 -960 418426 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 421626 -960 421738 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 428250 -960 428362 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 431562 -960 431674 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 163290 -960 163402 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 434874 -960 434986 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 438186 -960 438298 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 444810 -960 444922 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 448122 -960 448234 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 451434 -960 451546 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 454746 -960 454858 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 461370 -960 461482 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 464682 -960 464794 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 166602 -960 166714 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 137898 -960 138010 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 469098 -960 469210 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 472410 -960 472522 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 479034 -960 479146 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 482346 -960 482458 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 485658 -960 485770 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 488970 -960 489082 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 495594 -960 495706 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 498906 -960 499018 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 171018 -960 171130 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 502218 -960 502330 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 505530 -960 505642 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 512154 -960 512266 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 515466 -960 515578 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 518778 -960 518890 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 522090 -960 522202 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 528714 -960 528826 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 532026 -960 532138 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 174330 -960 174442 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 535338 -960 535450 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 538650 -960 538762 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 545274 -960 545386 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 548586 -960 548698 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 551898 -960 552010 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 555210 -960 555322 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 177642 -960 177754 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 180954 -960 181066 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 184266 -960 184378 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 187578 -960 187690 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 190890 -960 191002 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 194202 -960 194314 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 197514 -960 197626 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 200826 -960 200938 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 204138 -960 204250 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 207450 -960 207562 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 210762 -960 210874 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 214074 -960 214186 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 217386 -960 217498 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 220698 -960 220810 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 224010 -960 224122 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 227322 -960 227434 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 230634 -960 230746 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 233946 -960 234058 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 144522 -960 144634 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 237258 -960 237370 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 240570 -960 240682 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 243882 -960 243994 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 247194 -960 247306 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 250506 -960 250618 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 253818 -960 253930 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 257130 -960 257242 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 260442 -960 260554 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 263754 -960 263866 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 267066 -960 267178 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 147834 -960 147946 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 270378 -960 270490 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 273690 -960 273802 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 277002 -960 277114 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 280314 -960 280426 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283626 -960 283738 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286938 -960 287050 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290250 -960 290362 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293562 -960 293674 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 296874 -960 296986 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300186 -960 300298 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 151146 -960 151258 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 303498 -960 303610 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 306810 -960 306922 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 310122 -960 310234 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 313434 -960 313546 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 316746 -960 316858 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 320058 -960 320170 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 323370 -960 323482 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 326682 -960 326794 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 329994 -960 330106 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 333306 -960 333418 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 154458 -960 154570 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 336618 -960 336730 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 339930 -960 340042 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 343242 -960 343354 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 346554 -960 346666 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 349866 -960 349978 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 353178 -960 353290 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 356490 -960 356602 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 359802 -960 359914 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 363114 -960 363226 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 366426 -960 366538 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 369738 -960 369850 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 373050 -960 373162 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 376362 -960 376474 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 379674 -960 379786 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 382986 -960 383098 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 386298 -960 386410 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 389610 -960 389722 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 392922 -960 393034 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 396234 -960 396346 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 399546 -960 399658 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 161082 -960 161194 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 402858 -960 402970 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 406170 -960 406282 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 409482 -960 409594 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 412794 -960 412906 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 416106 -960 416218 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 419418 -960 419530 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 422730 -960 422842 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 426042 -960 426154 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 429354 -960 429466 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 432666 -960 432778 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 164394 -960 164506 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 435978 -960 436090 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 439290 -960 439402 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 445914 -960 446026 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 449226 -960 449338 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 452538 -960 452650 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 455850 -960 455962 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 462474 -960 462586 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 465786 -960 465898 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 167706 -960 167818 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 139002 -960 139114 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 470202 -960 470314 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 473514 -960 473626 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 476826 -960 476938 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 480138 -960 480250 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 483450 -960 483562 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 486762 -960 486874 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 490074 -960 490186 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 493386 -960 493498 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 496698 -960 496810 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 500010 -960 500122 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 172122 -960 172234 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 503322 -960 503434 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 506634 -960 506746 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 509946 -960 510058 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 513258 -960 513370 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 516570 -960 516682 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 519882 -960 519994 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 523194 -960 523306 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 526506 -960 526618 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 529818 -960 529930 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 533130 -960 533242 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 536442 -960 536554 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 539754 -960 539866 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 543066 -960 543178 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 546378 -960 546490 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 549690 -960 549802 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 553002 -960 553114 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 556314 -960 556426 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 559626 -960 559738 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 178746 -960 178858 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 182058 -960 182170 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 185370 -960 185482 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 188682 -960 188794 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 195306 -960 195418 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 198618 -960 198730 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 201930 -960 202042 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 142314 -960 142426 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 205242 -960 205354 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 211866 -960 211978 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 215178 -960 215290 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 218490 -960 218602 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 221802 -960 221914 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 228426 -960 228538 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 231738 -960 231850 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 235050 -960 235162 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 145626 -960 145738 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 238362 -960 238474 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 244986 -960 245098 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 248298 -960 248410 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 251610 -960 251722 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 254922 -960 255034 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 261546 -960 261658 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 264858 -960 264970 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 268170 -960 268282 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 148938 -960 149050 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 271482 -960 271594 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 278106 -960 278218 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 281418 -960 281530 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284730 -960 284842 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 288042 -960 288154 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294666 -960 294778 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 297978 -960 298090 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301290 -960 301402 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 152250 -960 152362 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 304602 -960 304714 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 311226 -960 311338 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 314538 -960 314650 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 317850 -960 317962 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 321162 -960 321274 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 324474 -960 324586 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 327786 -960 327898 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 331098 -960 331210 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 334410 -960 334522 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 155562 -960 155674 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 337722 -960 337834 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 341034 -960 341146 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 344346 -960 344458 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 347658 -960 347770 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 350970 -960 351082 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 354282 -960 354394 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 357594 -960 357706 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 360906 -960 361018 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 364218 -960 364330 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 367530 -960 367642 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 370842 -960 370954 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 374154 -960 374266 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 377466 -960 377578 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 380778 -960 380890 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 384090 -960 384202 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 387402 -960 387514 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 390714 -960 390826 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 394026 -960 394138 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 397338 -960 397450 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 400650 -960 400762 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 162186 -960 162298 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 403962 -960 404074 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 407274 -960 407386 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 410586 -960 410698 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 413898 -960 414010 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 417210 -960 417322 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 420522 -960 420634 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 423834 -960 423946 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 427146 -960 427258 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 430458 -960 430570 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 433770 -960 433882 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 165498 -960 165610 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 437082 -960 437194 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 440394 -960 440506 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 443706 -960 443818 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 447018 -960 447130 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 450330 -960 450442 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 453642 -960 453754 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 456954 -960 457066 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 460266 -960 460378 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 463578 -960 463690 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 466890 -960 467002 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 168810 -960 168922 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 560730 -960 560842 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 561834 -960 561946 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 562938 -960 563050 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 564042 -960 564154 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2316 -1244 -1696 705180 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2316 -1244 586240 -624 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2316 704560 586240 705180 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585620 -1244 586240 705180 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7964 2414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7964 38414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7964 74414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7964 110414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7964 146414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7964 182414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7964 218414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7964 254414 98000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 262000 254414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7964 290414 98000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 262000 290414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7964 326414 98000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 262000 326414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7964 362414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7964 398414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7964 434414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7964 470414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7964 506414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7964 542414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7964 578414 711900 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 2866 592960 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 38866 592960 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 74866 592960 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 110866 592960 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 146866 592960 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 182866 592960 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 218866 592960 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 254866 592960 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 290866 592960 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 326866 592960 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 362866 592960 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 398866 592960 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 434866 592960 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 470866 592960 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 506866 592960 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 542866 592960 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 578866 592960 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 614866 592960 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 650866 592960 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -9036 686866 592960 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -4236 -3164 -3616 707100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -4236 -3164 588160 -2544 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -4236 706480 588160 707100 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587540 -3164 588160 707100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7964 11414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7964 47414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7964 83414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7964 119414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7964 155414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7964 191414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7964 227414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7964 263414 98000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 262000 263414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7964 299414 98000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 262000 299414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7964 335414 98000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 262000 335414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7964 371414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7964 407414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7964 443414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7964 479414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7964 515414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7964 551414 711900 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 11866 592960 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 47866 592960 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 83866 592960 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 119866 592960 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 155866 592960 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 191866 592960 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 227866 592960 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 263866 592960 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 299866 592960 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 335866 592960 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 371866 592960 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 407866 592960 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 443866 592960 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 479866 592960 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 515866 592960 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 551866 592960 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 587866 592960 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 623866 592960 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 659866 592960 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -9036 695866 592960 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -6156 -5084 -5536 709020 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -6156 -5084 590080 -4464 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -6156 708400 590080 709020 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589460 -5084 590080 709020 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7964 20414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7964 56414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7964 92414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7964 128414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7964 164414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7964 200414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7964 236414 98000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 262000 236414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7964 272414 98000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 262000 272414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7964 308414 98000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 262000 308414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7964 344414 98000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 262000 344414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7964 380414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7964 416414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7964 452414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7964 488414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7964 524414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7964 560414 711900 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 20866 592960 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 56866 592960 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 92866 592960 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 128866 592960 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 164866 592960 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 200866 592960 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 236866 592960 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 272866 592960 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 308866 592960 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 344866 592960 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 380866 592960 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 416866 592960 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 452866 592960 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 488866 592960 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 524866 592960 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 560866 592960 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 596866 592960 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 632866 592960 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -9036 668866 592960 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -8076 -7004 -7456 710940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8076 -7004 592000 -6384 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8076 710320 592000 710940 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591380 -7004 592000 710940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7964 29414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7964 65414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7964 101414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7964 137414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7964 173414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7964 209414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7964 245414 98000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 262000 245414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7964 281414 98000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 262000 281414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7964 317414 98000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 262000 317414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7964 353414 98000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 262000 353414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7964 389414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7964 425414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7964 461414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7964 497414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7964 533414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7964 569414 711900 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 29866 592960 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 65866 592960 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 101866 592960 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 137866 592960 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 173866 592960 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 209866 592960 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 245866 592960 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 281866 592960 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 317866 592960 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 353866 592960 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 389866 592960 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 425866 592960 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 461866 592960 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 497866 592960 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 533866 592960 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 569866 592960 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 605866 592960 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 641866 592960 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -9036 677866 592960 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -7116 -6044 -6496 709980 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -7116 -6044 591040 -5424 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -7116 709360 591040 709980 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590420 -6044 591040 709980 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7964 24914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7964 60914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7964 96914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7964 132914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7964 168914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7964 204914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7964 240914 98000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 262000 240914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7964 276914 98000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 262000 276914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7964 312914 98000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 262000 312914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7964 348914 98000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 262000 348914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7964 384914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7964 420914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7964 456914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7964 492914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7964 528914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7964 564914 711900 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 25366 592960 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 61366 592960 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 97366 592960 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 133366 592960 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 169366 592960 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 205366 592960 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 241366 592960 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 277366 592960 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 313366 592960 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 349366 592960 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 385366 592960 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 421366 592960 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 457366 592960 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 493366 592960 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 529366 592960 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 565366 592960 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 601366 592960 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 637366 592960 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -9036 673366 592960 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -9036 -7964 -8416 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 -7964 592960 -7344 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 711280 592960 711900 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592340 -7964 592960 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7964 33914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7964 69914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7964 105914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7964 141914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7964 177914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7964 213914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7964 249914 98000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 262000 249914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7964 285914 98000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 262000 285914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7964 321914 98000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 262000 321914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7964 357914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7964 393914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7964 429914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7964 465914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7964 501914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7964 537914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7964 573914 711900 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 34366 592960 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 70366 592960 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 106366 592960 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 142366 592960 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 178366 592960 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 214366 592960 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 250366 592960 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 286366 592960 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 322366 592960 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 358366 592960 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 394366 592960 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 430366 592960 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 466366 592960 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 502366 592960 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 538366 592960 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 574366 592960 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 610366 592960 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 646366 592960 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -9036 682366 592960 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -3276 -2204 -2656 706140 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -3276 -2204 587200 -1584 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -3276 705520 587200 706140 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586580 -2204 587200 706140 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7964 6914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7964 42914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7964 78914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7964 114914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7964 150914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7964 186914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7964 222914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7964 258914 98000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 262000 258914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7964 294914 98000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 262000 294914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7964 330914 98000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 262000 330914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7964 366914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7964 402914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7964 438914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7964 474914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7964 510914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7964 546914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7964 582914 711900 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 7366 592960 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 43366 592960 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 79366 592960 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 115366 592960 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 151366 592960 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 187366 592960 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 223366 592960 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 259366 592960 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 295366 592960 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 331366 592960 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 367366 592960 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 403366 592960 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 439366 592960 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 475366 592960 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 511366 592960 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 547366 592960 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 583366 592960 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 619366 592960 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 655366 592960 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -9036 691366 592960 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -5196 -4124 -4576 708060 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -5196 -4124 589120 -3504 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -5196 707440 589120 708060 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588500 -4124 589120 708060 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7964 15914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7964 51914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7964 87914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7964 123914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7964 159914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7964 195914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7964 231914 98000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 262000 231914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7964 267914 98000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 262000 267914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7964 303914 98000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 262000 303914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7964 339914 98000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 262000 339914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7964 375914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7964 411914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7964 447914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7964 483914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7964 519914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7964 555914 711900 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 16366 592960 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 52366 592960 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 88366 592960 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 124366 592960 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 160366 592960 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 196366 592960 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 232366 592960 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 268366 592960 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 304366 592960 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 340366 592960 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 376366 592960 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 412366 592960 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 448366 592960 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 484366 592960 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 520366 592960 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 556366 592960 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 592366 592960 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 628366 592960 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 664366 592960 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -9036 700366 592960 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 19770 -960 19882 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 20874 -960 20986 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 21978 -960 22090 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 26394 -960 26506 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 63930 -960 64042 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 67242 -960 67354 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 70554 -960 70666 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 73866 -960 73978 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 77178 -960 77290 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 80490 -960 80602 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 83802 -960 83914 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 87114 -960 87226 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 90426 -960 90538 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 93738 -960 93850 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 30810 -960 30922 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 97050 -960 97162 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 100362 -960 100474 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 103674 -960 103786 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 106986 -960 107098 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 110298 -960 110410 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 113610 -960 113722 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 116922 -960 117034 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 120234 -960 120346 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 123546 -960 123658 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 126858 -960 126970 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 35226 -960 35338 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 130170 -960 130282 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 133482 -960 133594 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 39642 -960 39754 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 44058 -960 44170 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 47370 -960 47482 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 50682 -960 50794 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 53994 -960 54106 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 57306 -960 57418 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 60618 -960 60730 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 23082 -960 23194 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 27498 -960 27610 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 65034 -960 65146 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 68346 -960 68458 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 71658 -960 71770 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 78282 -960 78394 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 81594 -960 81706 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 84906 -960 85018 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 88218 -960 88330 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 94842 -960 94954 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 31914 -960 32026 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 98154 -960 98266 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 101466 -960 101578 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 104778 -960 104890 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 111402 -960 111514 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 114714 -960 114826 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 118026 -960 118138 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 121338 -960 121450 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 127962 -960 128074 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 36330 -960 36442 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 131274 -960 131386 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 134586 -960 134698 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 40746 -960 40858 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 45162 -960 45274 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 48474 -960 48586 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 51786 -960 51898 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 55098 -960 55210 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 61722 -960 61834 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 28602 -960 28714 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 66138 -960 66250 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 69450 -960 69562 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 72762 -960 72874 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 76074 -960 76186 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 79386 -960 79498 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 82698 -960 82810 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 86010 -960 86122 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 89322 -960 89434 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 92634 -960 92746 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 95946 -960 96058 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 33018 -960 33130 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 99258 -960 99370 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 102570 -960 102682 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 105882 -960 105994 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 109194 -960 109306 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 112506 -960 112618 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 115818 -960 115930 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 119130 -960 119242 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 122442 -960 122554 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 125754 -960 125866 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 129066 -960 129178 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 37434 -960 37546 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 132378 -960 132490 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 135690 -960 135802 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 46266 -960 46378 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 49578 -960 49690 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 52890 -960 53002 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 56202 -960 56314 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 59514 -960 59626 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 62826 -960 62938 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 29706 -960 29818 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 34122 -960 34234 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 38538 -960 38650 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 42954 -960 43066 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
