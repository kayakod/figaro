magic
tech sky130A
magscale 1 2
timestamp 1654675377
<< obsli1 >>
rect 1104 2159 118864 157777
<< obsm1 >>
rect 106 2128 119862 157808
<< metal2 >>
rect 2226 159200 2282 160000
rect 6642 159200 6698 160000
rect 11058 159200 11114 160000
rect 15474 159200 15530 160000
rect 19982 159200 20038 160000
rect 24398 159200 24454 160000
rect 28814 159200 28870 160000
rect 33322 159200 33378 160000
rect 37738 159200 37794 160000
rect 42154 159200 42210 160000
rect 46570 159200 46626 160000
rect 51078 159200 51134 160000
rect 55494 159200 55550 160000
rect 59910 159200 59966 160000
rect 64418 159200 64474 160000
rect 68834 159200 68890 160000
rect 73250 159200 73306 160000
rect 77758 159200 77814 160000
rect 82174 159200 82230 160000
rect 86590 159200 86646 160000
rect 91006 159200 91062 160000
rect 95514 159200 95570 160000
rect 99930 159200 99986 160000
rect 104346 159200 104402 160000
rect 108854 159200 108910 160000
rect 113270 159200 113326 160000
rect 117686 159200 117742 160000
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57978 0 58034 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60646 0 60702 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68650 0 68706 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78218 0 78274 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80610 0 80666 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81346 0 81402 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83554 0 83610 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87418 0 87474 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89626 0 89682 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92018 0 92074 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93306 0 93362 800
rect 93490 0 93546 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94502 0 94558 800
rect 94686 0 94742 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 95974 0 96030 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97906 0 97962 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99562 0 99618 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100298 0 100354 800
rect 100574 0 100630 800
rect 100850 0 100906 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103518 0 103574 800
rect 103702 0 103758 800
rect 103978 0 104034 800
rect 104254 0 104310 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105174 0 105230 800
rect 105450 0 105506 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106370 0 106426 800
rect 106646 0 106702 800
rect 106922 0 106978 800
rect 107106 0 107162 800
rect 107382 0 107438 800
rect 107658 0 107714 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108394 0 108450 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109038 0 109094 800
rect 109314 0 109370 800
rect 109590 0 109646 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110510 0 110566 800
rect 110786 0 110842 800
rect 111062 0 111118 800
rect 111246 0 111302 800
rect 111522 0 111578 800
rect 111798 0 111854 800
rect 111982 0 112038 800
rect 112258 0 112314 800
rect 112534 0 112590 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113178 0 113234 800
rect 113454 0 113510 800
rect 113730 0 113786 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115202 0 115258 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 115938 0 115994 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117318 0 117374 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118054 0 118110 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119526 0 119582 800
rect 119802 0 119858 800
<< obsm2 >>
rect 112 159144 2170 159338
rect 2338 159144 6586 159338
rect 6754 159144 11002 159338
rect 11170 159144 15418 159338
rect 15586 159144 19926 159338
rect 20094 159144 24342 159338
rect 24510 159144 28758 159338
rect 28926 159144 33266 159338
rect 33434 159144 37682 159338
rect 37850 159144 42098 159338
rect 42266 159144 46514 159338
rect 46682 159144 51022 159338
rect 51190 159144 55438 159338
rect 55606 159144 59854 159338
rect 60022 159144 64362 159338
rect 64530 159144 68778 159338
rect 68946 159144 73194 159338
rect 73362 159144 77702 159338
rect 77870 159144 82118 159338
rect 82286 159144 86534 159338
rect 86702 159144 90950 159338
rect 91118 159144 95458 159338
rect 95626 159144 99874 159338
rect 100042 159144 104290 159338
rect 104458 159144 108798 159338
rect 108966 159144 113214 159338
rect 113382 159144 117630 159338
rect 117798 159144 119856 159338
rect 112 856 119856 159144
rect 222 800 238 856
rect 406 800 514 856
rect 682 800 698 856
rect 866 800 974 856
rect 1142 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1710 856
rect 1878 800 1986 856
rect 2154 800 2170 856
rect 2338 800 2446 856
rect 2614 800 2722 856
rect 2890 800 2906 856
rect 3074 800 3182 856
rect 3350 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3918 856
rect 4086 800 4102 856
rect 4270 800 4378 856
rect 4546 800 4654 856
rect 4822 800 4838 856
rect 5006 800 5114 856
rect 5282 800 5390 856
rect 5558 800 5574 856
rect 5742 800 5850 856
rect 6018 800 6126 856
rect 6294 800 6310 856
rect 6478 800 6586 856
rect 6754 800 6862 856
rect 7030 800 7046 856
rect 7214 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7782 856
rect 7950 800 8058 856
rect 8226 800 8242 856
rect 8410 800 8518 856
rect 8686 800 8794 856
rect 8962 800 8978 856
rect 9146 800 9254 856
rect 9422 800 9530 856
rect 9698 800 9714 856
rect 9882 800 9990 856
rect 10158 800 10266 856
rect 10434 800 10450 856
rect 10618 800 10726 856
rect 10894 800 11002 856
rect 11170 800 11186 856
rect 11354 800 11462 856
rect 11630 800 11646 856
rect 11814 800 11922 856
rect 12090 800 12198 856
rect 12366 800 12382 856
rect 12550 800 12658 856
rect 12826 800 12934 856
rect 13102 800 13118 856
rect 13286 800 13394 856
rect 13562 800 13670 856
rect 13838 800 13854 856
rect 14022 800 14130 856
rect 14298 800 14406 856
rect 14574 800 14590 856
rect 14758 800 14866 856
rect 15034 800 15050 856
rect 15218 800 15326 856
rect 15494 800 15602 856
rect 15770 800 15786 856
rect 15954 800 16062 856
rect 16230 800 16338 856
rect 16506 800 16522 856
rect 16690 800 16798 856
rect 16966 800 17074 856
rect 17242 800 17258 856
rect 17426 800 17534 856
rect 17702 800 17810 856
rect 17978 800 17994 856
rect 18162 800 18270 856
rect 18438 800 18546 856
rect 18714 800 18730 856
rect 18898 800 19006 856
rect 19174 800 19190 856
rect 19358 800 19466 856
rect 19634 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20478 856
rect 20646 800 20662 856
rect 20830 800 20938 856
rect 21106 800 21214 856
rect 21382 800 21398 856
rect 21566 800 21674 856
rect 21842 800 21950 856
rect 22118 800 22134 856
rect 22302 800 22410 856
rect 22578 800 22594 856
rect 22762 800 22870 856
rect 23038 800 23146 856
rect 23314 800 23330 856
rect 23498 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24066 856
rect 24234 800 24342 856
rect 24510 800 24618 856
rect 24786 800 24802 856
rect 24970 800 25078 856
rect 25246 800 25354 856
rect 25522 800 25538 856
rect 25706 800 25814 856
rect 25982 800 26090 856
rect 26258 800 26274 856
rect 26442 800 26550 856
rect 26718 800 26734 856
rect 26902 800 27010 856
rect 27178 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27746 856
rect 27914 800 28022 856
rect 28190 800 28206 856
rect 28374 800 28482 856
rect 28650 800 28758 856
rect 28926 800 28942 856
rect 29110 800 29218 856
rect 29386 800 29494 856
rect 29662 800 29678 856
rect 29846 800 29954 856
rect 30122 800 30138 856
rect 30306 800 30414 856
rect 30582 800 30690 856
rect 30858 800 30874 856
rect 31042 800 31150 856
rect 31318 800 31426 856
rect 31594 800 31610 856
rect 31778 800 31886 856
rect 32054 800 32162 856
rect 32330 800 32346 856
rect 32514 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33082 856
rect 33250 800 33358 856
rect 33526 800 33634 856
rect 33802 800 33818 856
rect 33986 800 34094 856
rect 34262 800 34278 856
rect 34446 800 34554 856
rect 34722 800 34830 856
rect 34998 800 35014 856
rect 35182 800 35290 856
rect 35458 800 35566 856
rect 35734 800 35750 856
rect 35918 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36762 856
rect 36930 800 37038 856
rect 37206 800 37222 856
rect 37390 800 37498 856
rect 37666 800 37682 856
rect 37850 800 37958 856
rect 38126 800 38234 856
rect 38402 800 38418 856
rect 38586 800 38694 856
rect 38862 800 38970 856
rect 39138 800 39154 856
rect 39322 800 39430 856
rect 39598 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40442 856
rect 40610 800 40626 856
rect 40794 800 40902 856
rect 41070 800 41178 856
rect 41346 800 41362 856
rect 41530 800 41638 856
rect 41806 800 41822 856
rect 41990 800 42098 856
rect 42266 800 42374 856
rect 42542 800 42558 856
rect 42726 800 42834 856
rect 43002 800 43110 856
rect 43278 800 43294 856
rect 43462 800 43570 856
rect 43738 800 43846 856
rect 44014 800 44030 856
rect 44198 800 44306 856
rect 44474 800 44582 856
rect 44750 800 44766 856
rect 44934 800 45042 856
rect 45210 800 45226 856
rect 45394 800 45502 856
rect 45670 800 45778 856
rect 45946 800 45962 856
rect 46130 800 46238 856
rect 46406 800 46514 856
rect 46682 800 46698 856
rect 46866 800 46974 856
rect 47142 800 47250 856
rect 47418 800 47434 856
rect 47602 800 47710 856
rect 47878 800 47986 856
rect 48154 800 48170 856
rect 48338 800 48446 856
rect 48614 800 48722 856
rect 48890 800 48906 856
rect 49074 800 49182 856
rect 49350 800 49366 856
rect 49534 800 49642 856
rect 49810 800 49918 856
rect 50086 800 50102 856
rect 50270 800 50378 856
rect 50546 800 50654 856
rect 50822 800 50838 856
rect 51006 800 51114 856
rect 51282 800 51390 856
rect 51558 800 51574 856
rect 51742 800 51850 856
rect 52018 800 52126 856
rect 52294 800 52310 856
rect 52478 800 52586 856
rect 52754 800 52770 856
rect 52938 800 53046 856
rect 53214 800 53322 856
rect 53490 800 53506 856
rect 53674 800 53782 856
rect 53950 800 54058 856
rect 54226 800 54242 856
rect 54410 800 54518 856
rect 54686 800 54794 856
rect 54962 800 54978 856
rect 55146 800 55254 856
rect 55422 800 55530 856
rect 55698 800 55714 856
rect 55882 800 55990 856
rect 56158 800 56266 856
rect 56434 800 56450 856
rect 56618 800 56726 856
rect 56894 800 56910 856
rect 57078 800 57186 856
rect 57354 800 57462 856
rect 57630 800 57646 856
rect 57814 800 57922 856
rect 58090 800 58198 856
rect 58366 800 58382 856
rect 58550 800 58658 856
rect 58826 800 58934 856
rect 59102 800 59118 856
rect 59286 800 59394 856
rect 59562 800 59670 856
rect 59838 800 59854 856
rect 60022 800 60130 856
rect 60298 800 60314 856
rect 60482 800 60590 856
rect 60758 800 60866 856
rect 61034 800 61050 856
rect 61218 800 61326 856
rect 61494 800 61602 856
rect 61770 800 61786 856
rect 61954 800 62062 856
rect 62230 800 62338 856
rect 62506 800 62522 856
rect 62690 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63258 856
rect 63426 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63994 856
rect 64162 800 64270 856
rect 64438 800 64454 856
rect 64622 800 64730 856
rect 64898 800 65006 856
rect 65174 800 65190 856
rect 65358 800 65466 856
rect 65634 800 65742 856
rect 65910 800 65926 856
rect 66094 800 66202 856
rect 66370 800 66478 856
rect 66646 800 66662 856
rect 66830 800 66938 856
rect 67106 800 67214 856
rect 67382 800 67398 856
rect 67566 800 67674 856
rect 67842 800 67858 856
rect 68026 800 68134 856
rect 68302 800 68410 856
rect 68578 800 68594 856
rect 68762 800 68870 856
rect 69038 800 69146 856
rect 69314 800 69330 856
rect 69498 800 69606 856
rect 69774 800 69882 856
rect 70050 800 70066 856
rect 70234 800 70342 856
rect 70510 800 70618 856
rect 70786 800 70802 856
rect 70970 800 71078 856
rect 71246 800 71262 856
rect 71430 800 71538 856
rect 71706 800 71814 856
rect 71982 800 71998 856
rect 72166 800 72274 856
rect 72442 800 72550 856
rect 72718 800 72734 856
rect 72902 800 73010 856
rect 73178 800 73286 856
rect 73454 800 73470 856
rect 73638 800 73746 856
rect 73914 800 74022 856
rect 74190 800 74206 856
rect 74374 800 74482 856
rect 74650 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75218 856
rect 75386 800 75402 856
rect 75570 800 75678 856
rect 75846 800 75954 856
rect 76122 800 76138 856
rect 76306 800 76414 856
rect 76582 800 76690 856
rect 76858 800 76874 856
rect 77042 800 77150 856
rect 77318 800 77426 856
rect 77594 800 77610 856
rect 77778 800 77886 856
rect 78054 800 78162 856
rect 78330 800 78346 856
rect 78514 800 78622 856
rect 78790 800 78806 856
rect 78974 800 79082 856
rect 79250 800 79358 856
rect 79526 800 79542 856
rect 79710 800 79818 856
rect 79986 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80554 856
rect 80722 800 80830 856
rect 80998 800 81014 856
rect 81182 800 81290 856
rect 81458 800 81566 856
rect 81734 800 81750 856
rect 81918 800 82026 856
rect 82194 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82762 856
rect 82930 800 82946 856
rect 83114 800 83222 856
rect 83390 800 83498 856
rect 83666 800 83682 856
rect 83850 800 83958 856
rect 84126 800 84234 856
rect 84402 800 84418 856
rect 84586 800 84694 856
rect 84862 800 84970 856
rect 85138 800 85154 856
rect 85322 800 85430 856
rect 85598 800 85706 856
rect 85874 800 85890 856
rect 86058 800 86166 856
rect 86334 800 86350 856
rect 86518 800 86626 856
rect 86794 800 86902 856
rect 87070 800 87086 856
rect 87254 800 87362 856
rect 87530 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88098 856
rect 88266 800 88374 856
rect 88542 800 88558 856
rect 88726 800 88834 856
rect 89002 800 89110 856
rect 89278 800 89294 856
rect 89462 800 89570 856
rect 89738 800 89846 856
rect 90014 800 90030 856
rect 90198 800 90306 856
rect 90474 800 90490 856
rect 90658 800 90766 856
rect 90934 800 91042 856
rect 91210 800 91226 856
rect 91394 800 91502 856
rect 91670 800 91778 856
rect 91946 800 91962 856
rect 92130 800 92238 856
rect 92406 800 92514 856
rect 92682 800 92698 856
rect 92866 800 92974 856
rect 93142 800 93250 856
rect 93418 800 93434 856
rect 93602 800 93710 856
rect 93878 800 93894 856
rect 94062 800 94170 856
rect 94338 800 94446 856
rect 94614 800 94630 856
rect 94798 800 94906 856
rect 95074 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95642 856
rect 95810 800 95918 856
rect 96086 800 96102 856
rect 96270 800 96378 856
rect 96546 800 96654 856
rect 96822 800 96838 856
rect 97006 800 97114 856
rect 97282 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97850 856
rect 98018 800 98034 856
rect 98202 800 98310 856
rect 98478 800 98586 856
rect 98754 800 98770 856
rect 98938 800 99046 856
rect 99214 800 99322 856
rect 99490 800 99506 856
rect 99674 800 99782 856
rect 99950 800 100058 856
rect 100226 800 100242 856
rect 100410 800 100518 856
rect 100686 800 100794 856
rect 100962 800 100978 856
rect 101146 800 101254 856
rect 101422 800 101438 856
rect 101606 800 101714 856
rect 101882 800 101990 856
rect 102158 800 102174 856
rect 102342 800 102450 856
rect 102618 800 102726 856
rect 102894 800 102910 856
rect 103078 800 103186 856
rect 103354 800 103462 856
rect 103630 800 103646 856
rect 103814 800 103922 856
rect 104090 800 104198 856
rect 104366 800 104382 856
rect 104550 800 104658 856
rect 104826 800 104934 856
rect 105102 800 105118 856
rect 105286 800 105394 856
rect 105562 800 105578 856
rect 105746 800 105854 856
rect 106022 800 106130 856
rect 106298 800 106314 856
rect 106482 800 106590 856
rect 106758 800 106866 856
rect 107034 800 107050 856
rect 107218 800 107326 856
rect 107494 800 107602 856
rect 107770 800 107786 856
rect 107954 800 108062 856
rect 108230 800 108338 856
rect 108506 800 108522 856
rect 108690 800 108798 856
rect 108966 800 108982 856
rect 109150 800 109258 856
rect 109426 800 109534 856
rect 109702 800 109718 856
rect 109886 800 109994 856
rect 110162 800 110270 856
rect 110438 800 110454 856
rect 110622 800 110730 856
rect 110898 800 111006 856
rect 111174 800 111190 856
rect 111358 800 111466 856
rect 111634 800 111742 856
rect 111910 800 111926 856
rect 112094 800 112202 856
rect 112370 800 112478 856
rect 112646 800 112662 856
rect 112830 800 112938 856
rect 113106 800 113122 856
rect 113290 800 113398 856
rect 113566 800 113674 856
rect 113842 800 113858 856
rect 114026 800 114134 856
rect 114302 800 114410 856
rect 114578 800 114594 856
rect 114762 800 114870 856
rect 115038 800 115146 856
rect 115314 800 115330 856
rect 115498 800 115606 856
rect 115774 800 115882 856
rect 116050 800 116066 856
rect 116234 800 116342 856
rect 116510 800 116526 856
rect 116694 800 116802 856
rect 116970 800 117078 856
rect 117246 800 117262 856
rect 117430 800 117538 856
rect 117706 800 117814 856
rect 117982 800 117998 856
rect 118166 800 118274 856
rect 118442 800 118550 856
rect 118718 800 118734 856
rect 118902 800 119010 856
rect 119178 800 119286 856
rect 119454 800 119470 856
rect 119638 800 119746 856
<< metal3 >>
rect 0 158040 800 158160
rect 119200 158040 120000 158160
rect 119200 154504 120000 154624
rect 0 154232 800 154352
rect 119200 150968 120000 151088
rect 0 150424 800 150544
rect 119200 147432 120000 147552
rect 0 146616 800 146736
rect 119200 143896 120000 144016
rect 0 142808 800 142928
rect 119200 140360 120000 140480
rect 0 139000 800 139120
rect 119200 136824 120000 136944
rect 0 135192 800 135312
rect 119200 133152 120000 133272
rect 0 131384 800 131504
rect 119200 129616 120000 129736
rect 0 127576 800 127696
rect 119200 126080 120000 126200
rect 0 123768 800 123888
rect 119200 122544 120000 122664
rect 0 119960 800 120080
rect 119200 119008 120000 119128
rect 0 116152 800 116272
rect 119200 115472 120000 115592
rect 0 112344 800 112464
rect 119200 111936 120000 112056
rect 0 108536 800 108656
rect 119200 108400 120000 108520
rect 0 104728 800 104848
rect 119200 104728 120000 104848
rect 119200 101192 120000 101312
rect 0 100920 800 101040
rect 119200 97656 120000 97776
rect 0 97112 800 97232
rect 119200 94120 120000 94240
rect 0 93304 800 93424
rect 119200 90584 120000 90704
rect 0 89496 800 89616
rect 119200 87048 120000 87168
rect 0 85688 800 85808
rect 119200 83512 120000 83632
rect 0 81880 800 82000
rect 119200 79840 120000 79960
rect 0 78072 800 78192
rect 119200 76304 120000 76424
rect 0 74264 800 74384
rect 119200 72768 120000 72888
rect 0 70456 800 70576
rect 119200 69232 120000 69352
rect 0 66648 800 66768
rect 119200 65696 120000 65816
rect 0 62840 800 62960
rect 119200 62160 120000 62280
rect 0 59032 800 59152
rect 119200 58624 120000 58744
rect 0 55224 800 55344
rect 119200 55088 120000 55208
rect 0 51416 800 51536
rect 119200 51416 120000 51536
rect 119200 47880 120000 48000
rect 0 47608 800 47728
rect 119200 44344 120000 44464
rect 0 43800 800 43920
rect 119200 40808 120000 40928
rect 0 39992 800 40112
rect 119200 37272 120000 37392
rect 0 36184 800 36304
rect 119200 33736 120000 33856
rect 0 32376 800 32496
rect 119200 30200 120000 30320
rect 0 28568 800 28688
rect 119200 26528 120000 26648
rect 0 24760 800 24880
rect 119200 22992 120000 23112
rect 0 20952 800 21072
rect 119200 19456 120000 19576
rect 0 17144 800 17264
rect 119200 15920 120000 16040
rect 0 13336 800 13456
rect 119200 12384 120000 12504
rect 0 9528 800 9648
rect 119200 8848 120000 8968
rect 0 5720 800 5840
rect 119200 5312 120000 5432
rect 0 1912 800 2032
rect 119200 1776 120000 1896
<< obsm3 >>
rect 880 157960 119120 158133
rect 800 154704 119200 157960
rect 800 154432 119120 154704
rect 880 154424 119120 154432
rect 880 154152 119200 154424
rect 800 151168 119200 154152
rect 800 150888 119120 151168
rect 800 150624 119200 150888
rect 880 150344 119200 150624
rect 800 147632 119200 150344
rect 800 147352 119120 147632
rect 800 146816 119200 147352
rect 880 146536 119200 146816
rect 800 144096 119200 146536
rect 800 143816 119120 144096
rect 800 143008 119200 143816
rect 880 142728 119200 143008
rect 800 140560 119200 142728
rect 800 140280 119120 140560
rect 800 139200 119200 140280
rect 880 138920 119200 139200
rect 800 137024 119200 138920
rect 800 136744 119120 137024
rect 800 135392 119200 136744
rect 880 135112 119200 135392
rect 800 133352 119200 135112
rect 800 133072 119120 133352
rect 800 131584 119200 133072
rect 880 131304 119200 131584
rect 800 129816 119200 131304
rect 800 129536 119120 129816
rect 800 127776 119200 129536
rect 880 127496 119200 127776
rect 800 126280 119200 127496
rect 800 126000 119120 126280
rect 800 123968 119200 126000
rect 880 123688 119200 123968
rect 800 122744 119200 123688
rect 800 122464 119120 122744
rect 800 120160 119200 122464
rect 880 119880 119200 120160
rect 800 119208 119200 119880
rect 800 118928 119120 119208
rect 800 116352 119200 118928
rect 880 116072 119200 116352
rect 800 115672 119200 116072
rect 800 115392 119120 115672
rect 800 112544 119200 115392
rect 880 112264 119200 112544
rect 800 112136 119200 112264
rect 800 111856 119120 112136
rect 800 108736 119200 111856
rect 880 108600 119200 108736
rect 880 108456 119120 108600
rect 800 108320 119120 108456
rect 800 104928 119200 108320
rect 880 104648 119120 104928
rect 800 101392 119200 104648
rect 800 101120 119120 101392
rect 880 101112 119120 101120
rect 880 100840 119200 101112
rect 800 97856 119200 100840
rect 800 97576 119120 97856
rect 800 97312 119200 97576
rect 880 97032 119200 97312
rect 800 94320 119200 97032
rect 800 94040 119120 94320
rect 800 93504 119200 94040
rect 880 93224 119200 93504
rect 800 90784 119200 93224
rect 800 90504 119120 90784
rect 800 89696 119200 90504
rect 880 89416 119200 89696
rect 800 87248 119200 89416
rect 800 86968 119120 87248
rect 800 85888 119200 86968
rect 880 85608 119200 85888
rect 800 83712 119200 85608
rect 800 83432 119120 83712
rect 800 82080 119200 83432
rect 880 81800 119200 82080
rect 800 80040 119200 81800
rect 800 79760 119120 80040
rect 800 78272 119200 79760
rect 880 77992 119200 78272
rect 800 76504 119200 77992
rect 800 76224 119120 76504
rect 800 74464 119200 76224
rect 880 74184 119200 74464
rect 800 72968 119200 74184
rect 800 72688 119120 72968
rect 800 70656 119200 72688
rect 880 70376 119200 70656
rect 800 69432 119200 70376
rect 800 69152 119120 69432
rect 800 66848 119200 69152
rect 880 66568 119200 66848
rect 800 65896 119200 66568
rect 800 65616 119120 65896
rect 800 63040 119200 65616
rect 880 62760 119200 63040
rect 800 62360 119200 62760
rect 800 62080 119120 62360
rect 800 59232 119200 62080
rect 880 58952 119200 59232
rect 800 58824 119200 58952
rect 800 58544 119120 58824
rect 800 55424 119200 58544
rect 880 55288 119200 55424
rect 880 55144 119120 55288
rect 800 55008 119120 55144
rect 800 51616 119200 55008
rect 880 51336 119120 51616
rect 800 48080 119200 51336
rect 800 47808 119120 48080
rect 880 47800 119120 47808
rect 880 47528 119200 47800
rect 800 44544 119200 47528
rect 800 44264 119120 44544
rect 800 44000 119200 44264
rect 880 43720 119200 44000
rect 800 41008 119200 43720
rect 800 40728 119120 41008
rect 800 40192 119200 40728
rect 880 39912 119200 40192
rect 800 37472 119200 39912
rect 800 37192 119120 37472
rect 800 36384 119200 37192
rect 880 36104 119200 36384
rect 800 33936 119200 36104
rect 800 33656 119120 33936
rect 800 32576 119200 33656
rect 880 32296 119200 32576
rect 800 30400 119200 32296
rect 800 30120 119120 30400
rect 800 28768 119200 30120
rect 880 28488 119200 28768
rect 800 26728 119200 28488
rect 800 26448 119120 26728
rect 800 24960 119200 26448
rect 880 24680 119200 24960
rect 800 23192 119200 24680
rect 800 22912 119120 23192
rect 800 21152 119200 22912
rect 880 20872 119200 21152
rect 800 19656 119200 20872
rect 800 19376 119120 19656
rect 800 17344 119200 19376
rect 880 17064 119200 17344
rect 800 16120 119200 17064
rect 800 15840 119120 16120
rect 800 13536 119200 15840
rect 880 13256 119200 13536
rect 800 12584 119200 13256
rect 800 12304 119120 12584
rect 800 9728 119200 12304
rect 880 9448 119200 9728
rect 800 9048 119200 9448
rect 800 8768 119120 9048
rect 800 5920 119200 8768
rect 880 5640 119200 5920
rect 800 5512 119200 5640
rect 800 5232 119120 5512
rect 800 2112 119200 5232
rect 880 1976 119200 2112
rect 880 1939 119120 1976
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
<< labels >>
rlabel metal3 s 119200 1776 120000 1896 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 119200 108400 120000 108520 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 119200 119008 120000 119128 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 119200 129616 120000 129736 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 119200 140360 120000 140480 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 119200 150968 120000 151088 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 117686 159200 117742 160000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 104346 159200 104402 160000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 91006 159200 91062 160000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 77758 159200 77814 160000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 64418 159200 64474 160000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 119200 12384 120000 12504 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 51078 159200 51134 160000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 37738 159200 37794 160000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 24398 159200 24454 160000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 11058 159200 11114 160000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 158040 800 158160 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 119200 22992 120000 23112 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 119200 33736 120000 33856 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 119200 44344 120000 44464 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 119200 55088 120000 55208 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 119200 65696 120000 65816 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 119200 76304 120000 76424 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 119200 87048 120000 87168 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 119200 97656 120000 97776 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 119200 8848 120000 8968 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 119200 115472 120000 115592 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 119200 126080 120000 126200 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 119200 136824 120000 136944 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 119200 147432 120000 147552 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 119200 158040 120000 158160 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 108854 159200 108910 160000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 95514 159200 95570 160000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82174 159200 82230 160000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 68834 159200 68890 160000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 55494 159200 55550 160000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 119200 19456 120000 19576 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 42154 159200 42210 160000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 28814 159200 28870 160000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 15474 159200 15530 160000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 2226 159200 2282 160000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 150424 800 150544 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 127576 800 127696 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 93304 800 93424 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 119200 30200 120000 30320 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 119200 40808 120000 40928 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 119200 51416 120000 51536 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 119200 62160 120000 62280 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 119200 72768 120000 72888 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 119200 83512 120000 83632 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 119200 94120 120000 94240 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 119200 104728 120000 104848 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 119200 5312 120000 5432 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 119200 111936 120000 112056 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 119200 122544 120000 122664 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 119200 133152 120000 133272 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 119200 143896 120000 144016 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 119200 154504 120000 154624 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 113270 159200 113326 160000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 99930 159200 99986 160000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 86590 159200 86646 160000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 73250 159200 73306 160000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 59910 159200 59966 160000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 119200 15920 120000 16040 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 46570 159200 46626 160000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 33322 159200 33378 160000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 19982 159200 20038 160000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 6642 159200 6698 160000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 154232 800 154352 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 119960 800 120080 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 119200 26528 120000 26648 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 119200 37272 120000 37392 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 119200 47880 120000 48000 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 119200 58624 120000 58744 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 119200 69232 120000 69352 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 119200 79840 120000 79960 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 119200 90584 120000 90704 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 119200 101192 120000 101312 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6367480
string GDS_FILE /home/kaya/Desktop/caravel_example/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/signoff/user_proj_example.magic.gds
string GDS_START 234958
<< end >>

